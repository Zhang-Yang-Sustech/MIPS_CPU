`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/01/05 19:55:32
// Design Name: 
// Module Name: Vga
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module vga_control(
input wire vga_clk,
input wire sys_rst,
input wire [11:0] pix_data,//��ĳ���������Ϣ
output reg [9:0] pix_x,
output reg [9:0] pix_y,
output wire[0:0] hsync,
output wire[0:0] vsync,
output reg [11:0] vga_rgb
);

parameter H_SYNC =10'd96; //��ͬ������
parameter H_BA=10'd48;
parameter H_VA = 10'd640; //�Ϸ���ʾ����
parameter H_TO=10'd800;

parameter V_SYNC =10'd2; //��ͬ������
parameter V_BA=10'd33;
parameter V_VA = 10'd480; //�Ϸ���ʾ����
parameter V_TO=10'd525;

reg[9:0] cnt_h=10'b00000_00001;
reg[9:0] cnt_v=10'b00000_00001;


    
        always@(posedge vga_clk,posedge sys_rst)begin
        if(sys_rst==1'b1)begin
            cnt_v<=10'b00000_00001;
            end
            else if( (cnt_h==H_TO)&& (cnt_v < V_TO  ) ) begin
                cnt_v<=cnt_v+10'b00000_00001;
            end
            else if( (cnt_h ==H_TO) &&(cnt_v == V_TO  )  ) begin
                cnt_v<=10'b00000_00001;
            end
            else begin
            cnt_v <=cnt_v;
            end
        end
        
        always@(posedge vga_clk,posedge sys_rst)begin
             if(sys_rst==1'b1)begin
       cnt_h<=0;
       end
       else if(cnt_h ==(H_TO) ) begin
           cnt_h<=10'b00000_00001;
       end
       else begin
       cnt_h<=cnt_h+10'b00000_00001;
       end
        end



           always@(posedge  vga_clk)begin
                  if( (cnt_h >=H_SYNC +H_BA-1'b1)&& (cnt_h <H_SYNC +H_BA + H_VA-1'b1) &&
                     (cnt_v >= V_SYNC +V_BA ) && (cnt_v <V_SYNC +V_BA + V_VA)  )begin
                        pix_x <=cnt_h -(H_SYNC +H_BA ) ;
                        pix_y <=cnt_v-(V_SYNC +V_BA );
                    end
                    else begin
                        pix_x<=10'b00000_00000;
                        pix_y<=10'b00000_00000;
                    end
            end
            
                always@(posedge  vga_clk)begin
                          if( (cnt_h >=H_SYNC +H_BA)&& (cnt_h <H_SYNC +H_BA + H_VA) &&
                             (cnt_v >= V_SYNC +V_BA ) && (cnt_v <V_SYNC +V_BA + V_VA)  )begin
                              vga_rgb<=pix_data;
                            end
                            else begin
                                vga_rgb<=12'b0000_0000_0000;
                            end
                    end
            
            assign hsync =(cnt_h <=H_SYNC  ? 1'b0:1'b1);
            assign vsync =(cnt_v <= V_SYNC  ? 1'b0 :1'b1);
            
 endmodule

module vga_draw(//25MHz
input wire vga_clk,
input wire sys_rst,
input [31:0] a0,
input [31:0] a1,
input [31:0] a2,

input wire [9:0]pix_x,
input wire [9:0]pix_y,
output reg [11:0] pix_data
);
parameter off =4'b0000, no_st = 4'b0011, start = 4'b0111, movef = 4'b0110, moveb = 4'b0101;
//�ֶ�ģʽ���״̬���ֱ�Ϊ�ػ���δ�𲽡��𲽡�ǰ�������ˣ��ɿ������ҷ���
parameter wait_command=4'b1000,left_turning=4'b1001,right_turning=4'b1010,circle_turning=4'b1011,keep_go=4'b1110,semi_movef=4'b1111;
//�ֱ�Ϊ�ȴ�ָ���ת����ת����ͷ������ǰ�������ɿ������ҷ����ǰ��
parameter black = 12'h000, blue = 12'h00f, white = 12'hfff;

reg [255:0] char2 [63:0];//a0
reg [255:0] char3 [63:0];//a1
reg [255:0] char4 [63:0];//a2


reg [31:0] char22_0 [63:0];//��λ
reg [31:0] char22_1 [63:0];//ǧλ
reg [31:0] char22_2 [63:0];//��λ
reg [31:0] char22_3 [63:0];//ʮλ
reg [127:0] char22_4 [63:0];//��λ

reg [31:0] char33_0 [63:0];//��λ
reg [31:0] char33_1 [63:0];//ǧλ
reg [31:0] char33_2 [63:0];//��λ
reg [31:0] char33_3 [63:0];//ʮλ
reg [127:0] char33_4 [63:0];//��λ

reg [31:0] char44_0 [63:0];//��λ
reg [31:0] char44_1 [63:0];//ǧλ
reg [31:0] char44_2 [63:0];//��λ
reg [31:0] char44_3 [63:0];//ʮλ
reg [127:0] char44_4 [63:0];//��λ


reg [511:0] char   [479:0];//�ܵ����ؿ�
parameter w1 = 14'd10000, k1 = 10'd1000, h1 = 7'd100, t1 = 4'd10, o1 = 1'd1;


always@(posedge vga_clk) begin

char2[ 0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char2[ 1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char2[ 2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char2[ 3] <= 256'h0000000000000000000000000000000008000000000000000000000000000000;
char2[ 4] <= 256'h0000000000000000000000000000E0000E000000000000000000000000000000;
char2[ 5] <= 256'h0003C00000000000000000000000F0000F800000000000000000000000000000;
char2[ 6] <= 256'h0003C00000000000000000000000FC000F000000000000000000000000000000;
char2[ 7] <= 256'h0003C00000000000000000000000F0000E000000000000000000000000000000;
char2[ 8] <= 256'h0003C00000000000000000000001E0000E000000000000000000000000000000;
char2[ 9] <= 256'h0003C00000000000000000000001E0000E000400000000000000000000000000;
char2[10] <= 256'h000FFC0000000000000000000001C0000E000E00000000000000000000000000;
char2[11] <= 256'h003FFE00000000000007E0000003C0000E001F00000000000000000000000000;
char2[12] <= 256'h007FDF8000000000001FF8000003CFFFFFFFFF80000000000000000000000000;
char2[13] <= 256'h00F3CF8000000000003C1E00000387FFFFFFFFC0000000000000000000000000;
char2[14] <= 256'h01E3C7C00000000000700F00000782001E000000000000000000000000000000;
char2[15] <= 256'h03E3C7E00000000000E00700000700001E000000000000000000000000000000;
char2[16] <= 256'h03C3C7E00000000001E00380000F00001E000000000000000000000000000000;
char2[17] <= 256'h07C3C7E00000000003C003C0000E00001E000000000000000000000000000000;
char2[18] <= 256'h07C3CFE00000000003C001C0000E00001E000000000000000000000000000000;
char2[19] <= 256'h07C3CFE000000000078001E0001E00001E004000000000000000000000000000;
char2[20] <= 256'h07C3CFC000000000078000E0001C00601E00E000000000000000000000000000;
char2[21] <= 256'h07E3CFC000000000070000E0003F007FFFFFF800000000000000000000000000;
char2[22] <= 256'h07E3C000000000000F0000F0003F807FFFFFF800000000000000000000000000;
char2[23] <= 256'h07F3C000000000000F0000F0003F00780000F000000000000000000000000000;
char2[24] <= 256'h03FBC000000000000F0000F0007E00780000E000000000000000000000000000;
char2[25] <= 256'h03FFC000000000000F000070007E00780000E000000000000000000000000000;
char2[26] <= 256'h01FFC000000FF0001E00007800EE00780000E000000000000000000000000000;
char2[27] <= 256'h00FFC000007FFC001E00007800CE00780000E000000000000000000000000000;
char2[28] <= 256'h007FC00001F01E001E00007801CE00780000E000000000000000000000000000;
char2[29] <= 256'h003FE00003C00F001E000078018E00780000E000000000000000000000000000;
char2[30] <= 256'h001FF80003800F801E000078030E007FFFFFE000000000000000000000000000;
char2[31] <= 256'h000FFC00078007801E000078070E007FFFFFE000000000000000000000000000;
char2[32] <= 256'h0003FE00078007801E000078060E00780000E000001E00000000000000000000;
char2[33] <= 256'h0003FE00078007801E0000780C0E00780000E000007F80000000000000000000;
char2[34] <= 256'h0003FF00038007801E000078080E00780000E000007F80000000000000000000;
char2[35] <= 256'h0003FF80000007801E000078180E00780000E00000FF80000000000000000000;
char2[36] <= 256'h0003DFC000000F801E000078100E00780000E00000FFC0000000000000000000;
char2[37] <= 256'h0003CFC00003FF801E000078000E00780000E00000FF80000000000000000000;
char2[38] <= 256'h0003CFE0001FF7801E000078000E00780000E000007F80000000000000000000;
char2[39] <= 256'h0003C7E000FE07801E000078000E007FFFFFE000007F00000000000000000000;
char2[40] <= 256'h0003C3E001F007800F000070000E007FFFFFE000001C00000000000000000000;
char2[41] <= 256'h07C3C3E003C007800F0000F0000E00780000E000000000000000000000000000;
char2[42] <= 256'h0FE3C3E0078007800F0000F0000E00780000E000000000000000000000000000;
char2[43] <= 256'h0FE3C3E00F0007800F0000F0000E00780000E000000000000000000000000000;
char2[44] <= 256'h0FE3C3E00F000780070000E0000E00780000E000000000000000000000000000;
char2[45] <= 256'h0FE3C3E01E000780078001E0000E00780000E000000000000000000000000000;
char2[46] <= 256'h0FC3C3E01E000780078001E0000E00780000E000000000000000000000000000;
char2[47] <= 256'h0FC3C3E01E00078003C001C0000E00780000E000003E00000000000000000000;
char2[48] <= 256'h0FC3C3C01E00078403C003C0000E007FFFFFE000007F00000000000000000000;
char2[49] <= 256'h07C3C7C01E00078401E00380000E007FFFFFE00000FF80000000000000000000;
char2[50] <= 256'h03C3CF800F000F8400E00700000E00780000E00000FF80000000000000000000;
char2[51] <= 256'h01F3DF000F803F8400700F00000E00780000E00000FF80000000000000000000;
char2[52] <= 256'h00FFFC0007C0F788003C1E00000E00780000E00000FF80000000000000000000;
char2[53] <= 256'h003FF00003FFC3F8001FF800000E00780000E000007F80000000000000000000;
char2[54] <= 256'h0003C00000FF01E00007E000000E00780000E080007F00000000000000000000;
char2[55] <= 256'h0003C0000000000000000000000E00780000E1C0001C00000000000000000000;
char2[56] <= 256'h0003C0000000000000000000000E00780000E3E0000000000000000000000000;
char2[57] <= 256'h0003C0000000000000000000000EFFFFFFFFFFF0000000000000000000000000;
char2[58] <= 256'h0003C0000000000000000000000E7FFFFFFFFFF8000000000000000000000000;
char2[59] <= 256'h0003C0000000000000000000000E300000000000000000000000000000000000;
char2[60] <= 256'h0003C0000000000000000000000E000000000000000000000000000000000000;
char2[61] <= 256'h0000000000000000000000000008000000000000000000000000000000000000;
char2[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char2[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;/*C:\Users\86178\Desktop\???.BMP*/

char3[ 0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char3[ 1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char3[ 2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char3[ 3] <= 256'h0000000000000000000000000000000008000000000000000000000000000000;
char3[ 4] <= 256'h0000000000000000000000000000E0000E000000000000000000000000000000;
char3[ 5] <= 256'h0003C00000000000000000000000F0000F800000000000000000000000000000;
char3[ 6] <= 256'h0003C00000000000000000000000FC000F000000000000000000000000000000;
char3[ 7] <= 256'h0003C00000000000000000000000F0000E000000000000000000000000000000;
char3[ 8] <= 256'h0003C00000000000000000000001E0000E000000000000000000000000000000;
char3[ 9] <= 256'h0003C00000000000000000000001E0000E000400000000000000000000000000;
char3[10] <= 256'h000FFC0000000000000000000001C0000E000E00000000000000000000000000;
char3[11] <= 256'h003FFE0000000000000040000003C0000E001F00000000000000000000000000;
char3[12] <= 256'h007FDF80000000000000C0000003CFFFFFFFFF80000000000000000000000000;
char3[13] <= 256'h00F3CF80000000000001C000000387FFFFFFFFC0000000000000000000000000;
char3[14] <= 256'h01E3C7C0000000000007C000000782001E000000000000000000000000000000;
char3[15] <= 256'h03E3C7E00000000001FFC000000700001E000000000000000000000000000000;
char3[16] <= 256'h03C3C7E00000000001FFC000000F00001E000000000000000000000000000000;
char3[17] <= 256'h07C3C7E0000000000007C000000E00001E000000000000000000000000000000;
char3[18] <= 256'h07C3CFE0000000000003C000000E00001E000000000000000000000000000000;
char3[19] <= 256'h07C3CFE0000000000003C000001E00001E004000000000000000000000000000;
char3[20] <= 256'h07C3CFC0000000000003C000001C00601E00E000000000000000000000000000;
char3[21] <= 256'h07E3CFC0000000000003C000003F007FFFFFF800000000000000000000000000;
char3[22] <= 256'h07E3C000000000000003C000003F807FFFFFF800000000000000000000000000;
char3[23] <= 256'h07F3C000000000000003C000003F00780000F000000000000000000000000000;
char3[24] <= 256'h03FBC000000000000003C000007E00780000E000000000000000000000000000;
char3[25] <= 256'h03FFC000000000000003C000007E00780000E000000000000000000000000000;
char3[26] <= 256'h01FFC000000FF0000003C00000EE00780000E000000000000000000000000000;
char3[27] <= 256'h00FFC000007FFC000003C00000CE00780000E000000000000000000000000000;
char3[28] <= 256'h007FC00001F01E000003C00001CE00780000E000000000000000000000000000;
char3[29] <= 256'h003FE00003C00F000003C000018E00780000E000000000000000000000000000;
char3[30] <= 256'h001FF80003800F800003C000030E007FFFFFE000000000000000000000000000;
char3[31] <= 256'h000FFC00078007800003C000070E007FFFFFE000000000000000000000000000;
char3[32] <= 256'h0003FE00078007800003C000060E00780000E000001E00000000000000000000;
char3[33] <= 256'h0003FE00078007800003C0000C0E00780000E000007F80000000000000000000;
char3[34] <= 256'h0003FF00038007800003C000080E00780000E000007F80000000000000000000;
char3[35] <= 256'h0003FF80000007800003C000180E00780000E00000FF80000000000000000000;
char3[36] <= 256'h0003DFC000000F800003C000100E00780000E00000FFC0000000000000000000;
char3[37] <= 256'h0003CFC00003FF800003C000000E00780000E00000FF80000000000000000000;
char3[38] <= 256'h0003CFE0001FF7800003C000000E00780000E000007F80000000000000000000;
char3[39] <= 256'h0003C7E000FE07800003C000000E007FFFFFE000007F00000000000000000000;
char3[40] <= 256'h0003C3E001F007800003C000000E007FFFFFE000001C00000000000000000000;
char3[41] <= 256'h07C3C3E003C007800003C000000E00780000E000000000000000000000000000;
char3[42] <= 256'h0FE3C3E0078007800003C000000E00780000E000000000000000000000000000;
char3[43] <= 256'h0FE3C3E00F0007800003C000000E00780000E000000000000000000000000000;
char3[44] <= 256'h0FE3C3E00F0007800003C000000E00780000E000000000000000000000000000;
char3[45] <= 256'h0FE3C3E01E0007800003C000000E00780000E000000000000000000000000000;
char3[46] <= 256'h0FC3C3E01E0007800003C000000E00780000E000000000000000000000000000;
char3[47] <= 256'h0FC3C3E01E0007800003C000000E00780000E000003E00000000000000000000;
char3[48] <= 256'h0FC3C3C01E0007840003C000000E007FFFFFE000007F00000000000000000000;
char3[49] <= 256'h07C3C7C01E0007840003C000000E007FFFFFE00000FF80000000000000000000;
char3[50] <= 256'h03C3CF800F000F840003C000000E00780000E00000FF80000000000000000000;
char3[51] <= 256'h01F3DF000F803F840007E000000E00780000E00000FF80000000000000000000;
char3[52] <= 256'h00FFFC0007C0F788000FF000000E00780000E00000FF80000000000000000000;
char3[53] <= 256'h003FF00003FFC3F801FFFF80000E00780000E000007F80000000000000000000;
char3[54] <= 256'h0003C00000FF01E001FFFF80000E00780000E080007F00000000000000000000;
char3[55] <= 256'h0003C0000000000000000000000E00780000E1C0001C00000000000000000000;
char3[56] <= 256'h0003C0000000000000000000000E00780000E3E0000000000000000000000000;
char3[57] <= 256'h0003C0000000000000000000000EFFFFFFFFFFF0000000000000000000000000;
char3[58] <= 256'h0003C0000000000000000000000E7FFFFFFFFFF8000000000000000000000000;
char3[59] <= 256'h0003C0000000000000000000000E300000000000000000000000000000000000;
char3[60] <= 256'h0003C0000000000000000000000E000000000000000000000000000000000000;
char3[61] <= 256'h0000000000000000000000000008000000000000000000000000000000000000;
char3[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char3[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;/*C:\Users\86178\Desktop\???.BMP*/

char4[ 0] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char4[ 1] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char4[ 2] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char4[ 3] <= 256'h0000000000000000000000000000000008000000000000000000000000000000;
char4[ 4] <= 256'h0000000000000000000000000000E0000E000000000000000000000000000000;
char4[ 5] <= 256'h0003C00000000000000000000000F0000F800000000000000000000000000000;
char4[ 6] <= 256'h0003C00000000000000000000000FC000F000000000000000000000000000000;
char4[ 7] <= 256'h0003C00000000000000000000000F0000E000000000000000000000000000000;
char4[ 8] <= 256'h0003C00000000000000000000001E0000E000000000000000000000000000000;
char4[ 9] <= 256'h0003C00000000000000000000001E0000E000400000000000000000000000000;
char4[10] <= 256'h000FFC0000000000000000000001C0000E000E00000000000000000000000000;
char4[11] <= 256'h003FFE0000000000000FF0000003C0000E001F00000000000000000000000000;
char4[12] <= 256'h007FDF8000000000003FFE000003CFFFFFFFFF80000000000000000000000000;
char4[13] <= 256'h00F3CF800000000000F81F00000387FFFFFFFFC0000000000000000000000000;
char4[14] <= 256'h01E3C7C00000000001E00780000782001E000000000000000000000000000000;
char4[15] <= 256'h03E3C7E00000000003C003C0000700001E000000000000000000000000000000;
char4[16] <= 256'h03C3C7E000000000078001E0000F00001E000000000000000000000000000000;
char4[17] <= 256'h07C3C7E000000000070001E0000E00001E000000000000000000000000000000;
char4[18] <= 256'h07C3CFE000000000070000F0000E00001E000000000000000000000000000000;
char4[19] <= 256'h07C3CFE0000000000F0000F0001E00001E004000000000000000000000000000;
char4[20] <= 256'h07C3CFC0000000000F8000F0001C00601E00E000000000000000000000000000;
char4[21] <= 256'h07E3CFC0000000000F8000F0003F007FFFFFF800000000000000000000000000;
char4[22] <= 256'h07E3C000000000000FC000F0003F807FFFFFF800000000000000000000000000;
char4[23] <= 256'h07F3C000000000000FC000F0003F00780000F000000000000000000000000000;
char4[24] <= 256'h03FBC000000000000FC000F0007E00780000E000000000000000000000000000;
char4[25] <= 256'h03FFC00000000000078001E0007E00780000E000000000000000000000000000;
char4[26] <= 256'h01FFC000000FF000000001E000EE00780000E000000000000000000000000000;
char4[27] <= 256'h00FFC000007FFC00000001E000CE00780000E000000000000000000000000000;
char4[28] <= 256'h007FC00001F01E00000003C001CE00780000E000000000000000000000000000;
char4[29] <= 256'h003FE00003C00F00000003C0018E00780000E000000000000000000000000000;
char4[30] <= 256'h001FF80003800F8000000780030E007FFFFFE000000000000000000000000000;
char4[31] <= 256'h000FFC000780078000000F00070E007FFFFFE000000000000000000000000000;
char4[32] <= 256'h0003FE000780078000000E00060E00780000E000001E00000000000000000000;
char4[33] <= 256'h0003FE000780078000001C000C0E00780000E000007F80000000000000000000;
char4[34] <= 256'h0003FF000380078000003800080E00780000E000007F80000000000000000000;
char4[35] <= 256'h0003FF800000078000007000180E00780000E00000FF80000000000000000000;
char4[36] <= 256'h0003DFC000000F800000E000100E00780000E00000FFC0000000000000000000;
char4[37] <= 256'h0003CFC00003FF800001C000000E00780000E00000FF80000000000000000000;
char4[38] <= 256'h0003CFE0001FF78000038000000E00780000E000007F80000000000000000000;
char4[39] <= 256'h0003C7E000FE078000070000000E007FFFFFE000007F00000000000000000000;
char4[40] <= 256'h0003C3E001F00780000E0000000E007FFFFFE000001C00000000000000000000;
char4[41] <= 256'h07C3C3E003C00780001C0000000E00780000E000000000000000000000000000;
char4[42] <= 256'h0FE3C3E00780078000380000000E00780000E000000000000000000000000000;
char4[43] <= 256'h0FE3C3E00F00078000700000000E00780000E000000000000000000000000000;
char4[44] <= 256'h0FE3C3E00F00078000E00030000E00780000E000000000000000000000000000;
char4[45] <= 256'h0FE3C3E01E00078001C00030000E00780000E000000000000000000000000000;
char4[46] <= 256'h0FC3C3E01E00078003800030000E00780000E000000000000000000000000000;
char4[47] <= 256'h0FC3C3E01E00078007800030000E00780000E000003E00000000000000000000;
char4[48] <= 256'h0FC3C3C01E00078407000060000E007FFFFFE000007F00000000000000000000;
char4[49] <= 256'h07C3C7C01E0007840E0000E0000E007FFFFFE00000FF80000000000000000000;
char4[50] <= 256'h03C3CF800F000F841C0001E0000E00780000E00000FF80000000000000000000;
char4[51] <= 256'h01F3DF000F803F841FFFFFE0000E00780000E00000FF80000000000000000000;
char4[52] <= 256'h00FFFC0007C0F7881FFFFFE0000E00780000E00000FF80000000000000000000;
char4[53] <= 256'h003FF00003FFC3F81FFFFFE0000E00780000E000007F80000000000000000000;
char4[54] <= 256'h0003C00000FF01E01FFFFFE0000E00780000E080007F00000000000000000000;
char4[55] <= 256'h0003C0000000000000000000000E00780000E1C0001C00000000000000000000;
char4[56] <= 256'h0003C0000000000000000000000E00780000E3E0000000000000000000000000;
char4[57] <= 256'h0003C0000000000000000000000EFFFFFFFFFFF0000000000000000000000000;
char4[58] <= 256'h0003C0000000000000000000000E7FFFFFFFFFF8000000000000000000000000;
char4[59] <= 256'h0003C0000000000000000000000E300000000000000000000000000000000000;
char4[60] <= 256'h0003C0000000000000000000000E000000000000000000000000000000000000;
char4[61] <= 256'h0000000000000000000000000008000000000000000000000000000000000000;
char4[62] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;
char4[63] <= 256'h0000000000000000000000000000000000000000000000000000000000000000;/*C:\Users\86178\Desktop\???.BMP*/

 

           
         case(a0/w1)
                    4'd0: begin
                        char22_0[  0] <= 32'h00000000;
                        char22_0[  1] <= 32'h00000000;
                        char22_0[  2] <= 32'h00000000;
                        char22_0[  3] <= 32'h00000000;
                        char22_0[  4] <= 32'h00000000;
                        char22_0[  5] <= 32'h00000000;
                        char22_0[  6] <= 32'h00000000;
                        char22_0[  7] <= 32'h00000000;
                        char22_0[  8] <= 32'h00000000;
                        char22_0[  9] <= 32'h00000000;
                        char22_0[10] <= 32'h000FF000;
                        char22_0[11] <= 32'h003FFC00;
                        char22_0[12] <= 32'h007E7E00;
                        char22_0[13] <= 32'h00F81F00;
                        char22_0[14] <= 32'h01F00F80;
                        char22_0[15] <= 32'h03F00FC0;
                        char22_0[16] <= 32'h03E007C0;
                        char22_0[17] <= 32'h07E007E0;
                        char22_0[18] <= 32'h07C003E0;
                        char22_0[19] <= 32'h0FC003F0;
                        char22_0[20] <= 32'h0FC003F0;
                        char22_0[21] <= 32'h0FC003F0;
                        char22_0[22] <= 32'h1F8001F8;
                        char22_0[23] <= 32'h1F8001F8;
                        char22_0[24] <= 32'h1F8001F8;
                        char22_0[25] <= 32'h1F8001F8;
                        char22_0[26] <= 32'h1F8001F8;
                        char22_0[27] <= 32'h3F8001F8;
                        char22_0[28] <= 32'h3F8001F8;
                        char22_0[29] <= 32'h3F8001F8;
                        char22_0[30] <= 32'h3F8001F8;
                        char22_0[31] <= 32'h3F8001F8;
                        char22_0[32] <= 32'h3F8001F8;
                        char22_0[33] <= 32'h3F8001F8;
                        char22_0[34] <= 32'h3F8001F8;
                        char22_0[35] <= 32'h3F8001F8;
                        char22_0[36] <= 32'h3F8001F8;
                        char22_0[37] <= 32'h1F8001F8;
                        char22_0[38] <= 32'h1F8001F8;
                        char22_0[39] <= 32'h1F8001F8;
                        char22_0[40] <= 32'h1F8001F8;
                        char22_0[41] <= 32'h1F8001F0;
                        char22_0[42] <= 32'h0F8003F0;
                        char22_0[43] <= 32'h0FC003F0;
                        char22_0[44] <= 32'h0FC003F0;
                        char22_0[45] <= 32'h07C003E0;
                        char22_0[46] <= 32'h07E007E0;
                        char22_0[47] <= 32'h03E007C0;
                        char22_0[48] <= 32'h03F00FC0;
                        char22_0[49] <= 32'h01F00F80;
                        char22_0[50] <= 32'h00F81F00;
                        char22_0[51] <= 32'h007E7E00;
                        char22_0[52] <= 32'h003FFC00;
                        char22_0[53] <= 32'h000FF000;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//0
                    4'd1: begin
                        char22_0[  0] <= 32'h00000000;
                        char22_0[  1] <= 32'h00000000;
                        char22_0[  2] <= 32'h00000000;
                        char22_0[  3] <= 32'h00000000;
                        char22_0[  4] <= 32'h00000000;
                        char22_0[  5] <= 32'h00000000;
                        char22_0[  6] <= 32'h00000000;
                        char22_0[  7] <= 32'h00000000;
                        char22_0[  8] <= 32'h00000000;
                        char22_0[  9] <= 32'h00000000;
                        char22_0[10] <= 32'h0000E000;
                        char22_0[11] <= 32'h0001E000;
                        char22_0[12] <= 32'h0003E000;
                        char22_0[13] <= 32'h001FE000;
                        char22_0[14] <= 32'h03FFE000;
                        char22_0[15] <= 32'h03FFE000;
                        char22_0[16] <= 32'h0007E000;
                        char22_0[17] <= 32'h0007E000;
                        char22_0[18] <= 32'h0007E000;
                        char22_0[19] <= 32'h0007E000;
                        char22_0[20] <= 32'h0007E000;
                        char22_0[21] <= 32'h0007E000;
                        char22_0[22] <= 32'h0007E000;
                        char22_0[23] <= 32'h0007E000;
                        char22_0[24] <= 32'h0007E000;
                        char22_0[25] <= 32'h0007E000;
                        char22_0[26] <= 32'h0007E000;
                        char22_0[27] <= 32'h0007E000;
                        char22_0[28] <= 32'h0007E000;
                        char22_0[29] <= 32'h0007E000;
                        char22_0[30] <= 32'h0007E000;
                        char22_0[31] <= 32'h0007E000;
                        char22_0[32] <= 32'h0007E000;
                        char22_0[33] <= 32'h0007E000;
                        char22_0[34] <= 32'h0007E000;
                        char22_0[35] <= 32'h0007E000;
                        char22_0[36] <= 32'h0007E000;
                        char22_0[37] <= 32'h0007E000;
                        char22_0[38] <= 32'h0007E000;
                        char22_0[39] <= 32'h0007E000;
                        char22_0[40] <= 32'h0007E000;
                        char22_0[41] <= 32'h0007E000;
                        char22_0[42] <= 32'h0007E000;
                        char22_0[43] <= 32'h0007E000;
                        char22_0[44] <= 32'h0007E000;
                        char22_0[45] <= 32'h0007E000;
                        char22_0[46] <= 32'h0007E000;
                        char22_0[47] <= 32'h0007E000;
                        char22_0[48] <= 32'h0007E000;
                        char22_0[49] <= 32'h0007E000;
                        char22_0[50] <= 32'h0007E000;
                        char22_0[51] <= 32'h000FF800;
                        char22_0[52] <= 32'h03FFFFC0;
                        char22_0[53] <= 32'h03FFFFC0;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//1
                    4'd2: begin
                        char22_0[  0] <= 32'h00000000;
                        char22_0[  1] <= 32'h00000000;
                        char22_0[  2] <= 32'h00000000;
                        char22_0[  3] <= 32'h00000000;
                        char22_0[  4] <= 32'h00000000;
                        char22_0[  5] <= 32'h00000000;
                        char22_0[  6] <= 32'h00000000;
                        char22_0[  7] <= 32'h00000000;
                        char22_0[  8] <= 32'h00000000;
                        char22_0[  9] <= 32'h00000000;
                        char22_0[10] <= 32'h001FFC00;
                        char22_0[11] <= 32'h007FFF00;
                        char22_0[12] <= 32'h01F83F80;
                        char22_0[13] <= 32'h03E00FC0;
                        char22_0[14] <= 32'h07C007E0;
                        char22_0[15] <= 32'h078007E0;
                        char22_0[16] <= 32'h0F8003F0;
                        char22_0[17] <= 32'h0F8003F0;
                        char22_0[18] <= 32'h1F8003F0;
                        char22_0[19] <= 32'h1F8003F0;
                        char22_0[20] <= 32'h1FC003F0;
                        char22_0[21] <= 32'h1FC003F0;
                        char22_0[22] <= 32'h1FC003F0;
                        char22_0[23] <= 32'h0FC003F0;
                        char22_0[24] <= 32'h07C003F0;
                        char22_0[25] <= 32'h000003E0;
                        char22_0[26] <= 32'h000007E0;
                        char22_0[27] <= 32'h000007E0;
                        char22_0[28] <= 32'h00000FC0;
                        char22_0[29] <= 32'h00000F80;
                        char22_0[30] <= 32'h00001F80;
                        char22_0[31] <= 32'h00003F00;
                        char22_0[32] <= 32'h00003E00;
                        char22_0[33] <= 32'h00007C00;
                        char22_0[34] <= 32'h0000F800;
                        char22_0[35] <= 32'h0001F000;
                        char22_0[36] <= 32'h0003E000;
                        char22_0[37] <= 32'h0007C000;
                        char22_0[38] <= 32'h000F8000;
                        char22_0[39] <= 32'h001F0000;
                        char22_0[40] <= 32'h003E0000;
                        char22_0[41] <= 32'h007C0000;
                        char22_0[42] <= 32'h00F80000;
                        char22_0[43] <= 32'h01F00038;
                        char22_0[44] <= 32'h01E00038;
                        char22_0[45] <= 32'h03C00070;
                        char22_0[46] <= 32'h07800070;
                        char22_0[47] <= 32'h0F8000F0;
                        char22_0[48] <= 32'h0F0000F0;
                        char22_0[49] <= 32'h1E0003F0;
                        char22_0[50] <= 32'h3FFFFFF0;
                        char22_0[51] <= 32'h3FFFFFF0;
                        char22_0[52] <= 32'h3FFFFFE0;
                        char22_0[53] <= 32'h3FFFFFE0;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//2
                    4'd3: begin
                        char22_0[  0] <= 32'h00000000;
                        char22_0[  1] <= 32'h00000000;
                        char22_0[  2] <= 32'h00000000;
                        char22_0[  3] <= 32'h00000000;
                        char22_0[  4] <= 32'h00000000;
                        char22_0[  5] <= 32'h00000000;
                        char22_0[  6] <= 32'h00000000;
                        char22_0[  7] <= 32'h00000000;
                        char22_0[  8] <= 32'h00000000;
                        char22_0[  9] <= 32'h00000000;
                        char22_0[10] <= 32'h003FF000;
                        char22_0[11] <= 32'h00FFFC00;
                        char22_0[12] <= 32'h01F07E00;
                        char22_0[13] <= 32'h03C03F00;
                        char22_0[14] <= 32'h07801F80;
                        char22_0[15] <= 32'h0F800FC0;
                        char22_0[16] <= 32'h0F800FC0;
                        char22_0[17] <= 32'h0F8007E0;
                        char22_0[18] <= 32'h0FC007E0;
                        char22_0[19] <= 32'h0FC007E0;
                        char22_0[20] <= 32'h0FC007E0;
                        char22_0[21] <= 32'h07C007E0;
                        char22_0[22] <= 32'h000007E0;
                        char22_0[23] <= 32'h000007E0;
                        char22_0[24] <= 32'h000007C0;
                        char22_0[25] <= 32'h00000FC0;
                        char22_0[26] <= 32'h00000F80;
                        char22_0[27] <= 32'h00001F00;
                        char22_0[28] <= 32'h00007E00;
                        char22_0[29] <= 32'h0003FC00;
                        char22_0[30] <= 32'h001FF000;
                        char22_0[31] <= 32'h001FFC00;
                        char22_0[32] <= 32'h0000FF00;
                        char22_0[33] <= 32'h00001F80;
                        char22_0[34] <= 32'h00000FC0;
                        char22_0[35] <= 32'h000007E0;
                        char22_0[36] <= 32'h000003E0;
                        char22_0[37] <= 32'h000003F0;
                        char22_0[38] <= 32'h000003F0;
                        char22_0[39] <= 32'h000001F0;
                        char22_0[40] <= 32'h000001F8;
                        char22_0[41] <= 32'h000001F8;
                        char22_0[42] <= 32'h078001F8;
                        char22_0[43] <= 32'h0FC001F8;
                        char22_0[44] <= 32'h1FC001F8;
                        char22_0[45] <= 32'h1FC003F0;
                        char22_0[46] <= 32'h1FC003F0;
                        char22_0[47] <= 32'h1FC003E0;
                        char22_0[48] <= 32'h0F8007E0;
                        char22_0[49] <= 32'h0F8007C0;
                        char22_0[50] <= 32'h07C01F80;
                        char22_0[51] <= 32'h03F07F00;
                        char22_0[52] <= 32'h01FFFE00;
                        char22_0[53] <= 32'h003FF000;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//3
                    4'd4: begin
                        char22_0[  0] <= 32'h00000000;
                        char22_0[  1] <= 32'h00000000;
                        char22_0[  2] <= 32'h00000000;
                        char22_0[  3] <= 32'h00000000;
                        char22_0[  4] <= 32'h00000000;
                        char22_0[  5] <= 32'h00000000;
                        char22_0[  6] <= 32'h00000000;
                        char22_0[  7] <= 32'h00000000;
                        char22_0[  8] <= 32'h00000000;
                        char22_0[  9] <= 32'h00000000;
                        char22_0[10] <= 32'h00001F00;
                        char22_0[11] <= 32'h00001F00;
                        char22_0[12] <= 32'h00003F00;
                        char22_0[13] <= 32'h00003F00;
                        char22_0[14] <= 32'h00007F00;
                        char22_0[15] <= 32'h0000FF00;
                        char22_0[16] <= 32'h0000FF00;
                        char22_0[17] <= 32'h0001FF00;
                        char22_0[18] <= 32'h0003FF00;
                        char22_0[19] <= 32'h0003BF00;
                        char22_0[20] <= 32'h0007BF00;
                        char22_0[21] <= 32'h00073F00;
                        char22_0[22] <= 32'h000F3F00;
                        char22_0[23] <= 32'h001E3F00;
                        char22_0[24] <= 32'h001C3F00;
                        char22_0[25] <= 32'h003C3F00;
                        char22_0[26] <= 32'h00783F00;
                        char22_0[27] <= 32'h00783F00;
                        char22_0[28] <= 32'h00F03F00;
                        char22_0[29] <= 32'h00E03F00;
                        char22_0[30] <= 32'h01E03F00;
                        char22_0[31] <= 32'h03C03F00;
                        char22_0[32] <= 32'h03803F00;
                        char22_0[33] <= 32'h07803F00;
                        char22_0[34] <= 32'h0F003F00;
                        char22_0[35] <= 32'h0F003F00;
                        char22_0[36] <= 32'h1E003F00;
                        char22_0[37] <= 32'h1C003F00;
                        char22_0[38] <= 32'h3C003F00;
                        char22_0[39] <= 32'h7FFFFFFE;
                        char22_0[40] <= 32'h7FFFFFFE;
                        char22_0[41] <= 32'h00003F00;
                        char22_0[42] <= 32'h00003F00;
                        char22_0[43] <= 32'h00003F00;
                        char22_0[44] <= 32'h00003F00;
                        char22_0[45] <= 32'h00003F00;
                        char22_0[46] <= 32'h00003F00;
                        char22_0[47] <= 32'h00003F00;
                        char22_0[48] <= 32'h00003F00;
                        char22_0[49] <= 32'h00003F00;
                        char22_0[50] <= 32'h00003F00;
                        char22_0[51] <= 32'h00007F80;
                        char22_0[52] <= 32'h000FFFFC;
                        char22_0[53] <= 32'h000FFFFC;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//4
                    4'd5: begin
                        char22_0[  0] <= 32'h00000000;
                        char22_0[  1] <= 32'h00000000;
                        char22_0[  2] <= 32'h00000000;
                        char22_0[  3] <= 32'h00000000;
                        char22_0[  4] <= 32'h00000000;
                        char22_0[  5] <= 32'h00000000;
                        char22_0[  6] <= 32'h00000000;
                        char22_0[  7] <= 32'h00000000;
                        char22_0[  8] <= 32'h00000000;
                        char22_0[  9] <= 32'h00000000;
                        char22_0[10] <= 32'h00000000;
                        char22_0[11] <= 32'h03FFFFF0;
                        char22_0[12] <= 32'h03FFFFF0;
                        char22_0[13] <= 32'h03FFFFF0;
                        char22_0[14] <= 32'h03FFFFE0;
                        char22_0[15] <= 32'h03800000;
                        char22_0[16] <= 32'h03800000;
                        char22_0[17] <= 32'h03800000;
                        char22_0[18] <= 32'h03800000;
                        char22_0[19] <= 32'h03800000;
                        char22_0[20] <= 32'h07800000;
                        char22_0[21] <= 32'h07800000;
                        char22_0[22] <= 32'h07800000;
                        char22_0[23] <= 32'h07800000;
                        char22_0[24] <= 32'h07800000;
                        char22_0[25] <= 32'h07800000;
                        char22_0[26] <= 32'h078FF800;
                        char22_0[27] <= 32'h073FFE00;
                        char22_0[28] <= 32'h077FFF80;
                        char22_0[29] <= 32'h07FC3F80;
                        char22_0[30] <= 32'h07E00FC0;
                        char22_0[31] <= 32'h07C007E0;
                        char22_0[32] <= 32'h078007E0;
                        char22_0[33] <= 32'h078003F0;
                        char22_0[34] <= 32'h000003F0;
                        char22_0[35] <= 32'h000001F0;
                        char22_0[36] <= 32'h000001F8;
                        char22_0[37] <= 32'h000001F8;
                        char22_0[38] <= 32'h000001F8;
                        char22_0[39] <= 32'h000001F8;
                        char22_0[40] <= 32'h000001F8;
                        char22_0[41] <= 32'h078001F8;
                        char22_0[42] <= 32'h0FC001F8;
                        char22_0[43] <= 32'h1FC001F0;
                        char22_0[44] <= 32'h1FC001F0;
                        char22_0[45] <= 32'h1FC003F0;
                        char22_0[46] <= 32'h1F8003F0;
                        char22_0[47] <= 32'h1F8003E0;
                        char22_0[48] <= 32'h0F8007E0;
                        char22_0[49] <= 32'h078007C0;
                        char22_0[50] <= 32'h07C01F80;
                        char22_0[51] <= 32'h03F83F00;
                        char22_0[52] <= 32'h00FFFE00;
                        char22_0[53] <= 32'h003FF800;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//5
                    4'd6: begin
                        char22_0[0] <= 32'h00000000;
                        char22_0[1] <= 32'h00000000;
                        char22_0[2] <= 32'h00000000;
                        char22_0[3] <= 32'h00000000;
                        char22_0[4] <= 32'h00000000;
                        char22_0[5] <= 32'h00000000;
                        char22_0[6] <= 32'h00000000;
                        char22_0[7] <= 32'h00000000;
                        char22_0[8] <= 32'h00000000;
                        char22_0[9] <= 32'h00000000;
                        char22_0[10] <= 32'h0007FE00;
                        char22_0[11] <= 32'h001FFF80;
                        char22_0[12] <= 32'h003F0FC0;
                        char22_0[13] <= 32'h007C07C0;
                        char22_0[14] <= 32'h00F807E0;
                        char22_0[15] <= 32'h01F007E0;
                        char22_0[16] <= 32'h03E007E0;
                        char22_0[17] <= 32'h03C007E0;
                        char22_0[18] <= 32'h07C003C0;
                        char22_0[19] <= 32'h07C00000;
                        char22_0[20] <= 32'h0FC00000;
                        char22_0[21] <= 32'h0F800000;
                        char22_0[22] <= 32'h0F800000;
                        char22_0[23] <= 32'h1F800000;
                        char22_0[24] <= 32'h1F800000;
                        char22_0[25] <= 32'h1F800000;
                        char22_0[26] <= 32'h1F87FE00;
                        char22_0[27] <= 32'h1F9FFF80;
                        char22_0[28] <= 32'h1FBFFFC0;
                        char22_0[29] <= 32'h3FFE1FC0;
                        char22_0[30] <= 32'h3FF807E0;
                        char22_0[31] <= 32'h3FE003F0;
                        char22_0[32] <= 32'h3FE003F0;
                        char22_0[33] <= 32'h3FC001F8;
                        char22_0[34] <= 32'h3F8001F8;
                        char22_0[35] <= 32'h3F8001F8;
                        char22_0[36] <= 32'h3F8000F8;
                        char22_0[37] <= 32'h3F8000F8;
                        char22_0[38] <= 32'h3F8000F8;
                        char22_0[39] <= 32'h1F8000F8;
                        char22_0[40] <= 32'h1F8000F8;
                        char22_0[41] <= 32'h1F8000F8;
                        char22_0[42] <= 32'h1F8000F8;
                        char22_0[43] <= 32'h1F8000F8;
                        char22_0[44] <= 32'h0FC001F8;
                        char22_0[45] <= 32'h0FC001F8;
                        char22_0[46] <= 32'h0FC001F0;
                        char22_0[47] <= 32'h07E001F0;
                        char22_0[48] <= 32'h03E003E0;
                        char22_0[49] <= 32'h03F003E0;
                        char22_0[50] <= 32'h01F807C0;
                        char22_0[51] <= 32'h00FE1F80;
                        char22_0[52] <= 32'h007FFE00;
                        char22_0[53] <= 32'h001FF800;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//6
                    4'd7: begin
                        char22_0[0] <= 32'h00000000;
                        char22_0[1] <= 32'h00000000;
                        char22_0[2] <= 32'h00000000;
                        char22_0[3] <= 32'h00000000;
                        char22_0[4] <= 32'h00000000;
                        char22_0[5] <= 32'h00000000;
                        char22_0[6] <= 32'h00000000;
                        char22_0[7] <= 32'h00000000;
                        char22_0[8] <= 32'h00000000;
                        char22_0[9] <= 32'h00000000;
                        char22_0[10] <= 32'h00000000;
                        char22_0[11] <= 32'h07FFFFF8;
                        char22_0[12] <= 32'h07FFFFF8;
                        char22_0[13] <= 32'h07FFFFF8;
                        char22_0[14] <= 32'h0FFFFFF0;
                        char22_0[15] <= 32'h0FC000E0;
                        char22_0[16] <= 32'h0F8001E0;
                        char22_0[17] <= 32'h0F0001C0;
                        char22_0[18] <= 32'h0E0003C0;
                        char22_0[19] <= 32'h0E000780;
                        char22_0[20] <= 32'h1E000780;
                        char22_0[21] <= 32'h1C000F00;
                        char22_0[22] <= 32'h00000F00;
                        char22_0[23] <= 32'h00001E00;
                        char22_0[24] <= 32'h00001E00;
                        char22_0[25] <= 32'h00003C00;
                        char22_0[26] <= 32'h00003C00;
                        char22_0[27] <= 32'h00007800;
                        char22_0[28] <= 32'h00007800;
                        char22_0[29] <= 32'h0000F800;
                        char22_0[30] <= 32'h0000F000;
                        char22_0[31] <= 32'h0001F000;
                        char22_0[32] <= 32'h0001E000;
                        char22_0[33] <= 32'h0003E000;
                        char22_0[34] <= 32'h0003E000;
                        char22_0[35] <= 32'h0003E000;
                        char22_0[36] <= 32'h0007C000;
                        char22_0[37] <= 32'h0007C000;
                        char22_0[38] <= 32'h0007C000;
                        char22_0[39] <= 32'h000FC000;
                        char22_0[40] <= 32'h000FC000;
                        char22_0[41] <= 32'h000FC000;
                        char22_0[42] <= 32'h000FC000;
                        char22_0[43] <= 32'h001FC000;
                        char22_0[44] <= 32'h001FC000;
                        char22_0[45] <= 32'h001FC000;
                        char22_0[46] <= 32'h001FC000;
                        char22_0[47] <= 32'h001FC000;
                        char22_0[48] <= 32'h001FC000;
                        char22_0[49] <= 32'h001FC000;
                        char22_0[50] <= 32'h001FC000;
                        char22_0[51] <= 32'h001FC000;
                        char22_0[52] <= 32'h001FC000;
                        char22_0[53] <= 32'h000F8000;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//7
                    4'd8: begin
                        char22_0[0] <= 32'h00000000;
                        char22_0[1] <= 32'h00000000;
                        char22_0[2] <= 32'h00000000;
                        char22_0[3] <= 32'h00000000;
                        char22_0[4] <= 32'h00000000;
                        char22_0[5] <= 32'h00000000;
                        char22_0[6] <= 32'h00000000;
                        char22_0[7] <= 32'h00000000;
                        char22_0[8] <= 32'h00000000;
                        char22_0[9] <= 32'h00000000;
                        char22_0[10] <= 32'h003FF800;
                        char22_0[11] <= 32'h00FFFE00;
                        char22_0[12] <= 32'h01F81F80;
                        char22_0[13] <= 32'h03E00FC0;
                        char22_0[14] <= 32'h07C003E0;
                        char22_0[15] <= 32'h0F8003E0;
                        char22_0[16] <= 32'h0F8001F0;
                        char22_0[17] <= 32'h1F0001F0;
                        char22_0[18] <= 32'h1F0001F0;
                        char22_0[19] <= 32'h1F0001F0;
                        char22_0[20] <= 32'h1F0001F0;
                        char22_0[21] <= 32'h1F0001F0;
                        char22_0[22] <= 32'h1F8001F0;
                        char22_0[23] <= 32'h1FC001F0;
                        char22_0[24] <= 32'h0FC001F0;
                        char22_0[25] <= 32'h0FF003E0;
                        char22_0[26] <= 32'h07F803C0;
                        char22_0[27] <= 32'h03FE0F80;
                        char22_0[28] <= 32'h01FF9F00;
                        char22_0[29] <= 32'h00FFFE00;
                        char22_0[30] <= 32'h003FF800;
                        char22_0[31] <= 32'h007FFC00;
                        char22_0[32] <= 32'h01F7FF00;
                        char22_0[33] <= 32'h03E1FF80;
                        char22_0[34] <= 32'h07C07FC0;
                        char22_0[35] <= 32'h0F801FE0;
                        char22_0[36] <= 32'h0F800FE0;
                        char22_0[37] <= 32'h1F0007F0;
                        char22_0[38] <= 32'h1F0003F0;
                        char22_0[39] <= 32'h3E0001F8;
                        char22_0[40] <= 32'h3E0001F8;
                        char22_0[41] <= 32'h3E0001F8;
                        char22_0[42] <= 32'h3E0000F8;
                        char22_0[43] <= 32'h3E0000F8;
                        char22_0[44] <= 32'h3E0000F8;
                        char22_0[45] <= 32'h3E0000F8;
                        char22_0[46] <= 32'h1F0001F0;
                        char22_0[47] <= 32'h1F0001F0;
                        char22_0[48] <= 32'h0F8003E0;
                        char22_0[49] <= 32'h0FC003E0;
                        char22_0[50] <= 32'h07E007C0;
                        char22_0[51] <= 32'h01F83F80;
                        char22_0[52] <= 32'h00FFFE00;
                        char22_0[53] <= 32'h003FF800;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//8
                    4'd9: begin
                        char22_0[0] <= 32'h00000000;
                        char22_0[1] <= 32'h00000000;
                        char22_0[2] <= 32'h00000000;
                        char22_0[3] <= 32'h00000000;
                        char22_0[4] <= 32'h00000000;
                        char22_0[5] <= 32'h00000000;
                        char22_0[6] <= 32'h00000000;
                        char22_0[7] <= 32'h00000000;
                        char22_0[8] <= 32'h00000000;
                        char22_0[9] <= 32'h00000000;
                        char22_0[10] <= 32'h003FF000;
                        char22_0[11] <= 32'h00FFFC00;
                        char22_0[12] <= 32'h01F83F00;
                        char22_0[13] <= 32'h03E01F80;
                        char22_0[14] <= 32'h07C00F80;
                        char22_0[15] <= 32'h0FC007C0;
                        char22_0[16] <= 32'h0F8003E0;
                        char22_0[17] <= 32'h1F8003E0;
                        char22_0[18] <= 32'h1F0003F0;
                        char22_0[19] <= 32'h1F0003F0;
                        char22_0[20] <= 32'h3F0001F0;
                        char22_0[21] <= 32'h3F0001F0;
                        char22_0[22] <= 32'h3F0001F8;
                        char22_0[23] <= 32'h3F0001F8;
                        char22_0[24] <= 32'h3F0001F8;
                        char22_0[25] <= 32'h3F0001F8;
                        char22_0[26] <= 32'h3F0001F8;
                        char22_0[27] <= 32'h3F0001F8;
                        char22_0[28] <= 32'h3F0003F8;
                        char22_0[29] <= 32'h1F8003F8;
                        char22_0[30] <= 32'h1F8007F8;
                        char22_0[31] <= 32'h1F800FF8;
                        char22_0[32] <= 32'h0FC01FF8;
                        char22_0[33] <= 32'h0FE03FF8;
                        char22_0[34] <= 32'h07F8FDF8;
                        char22_0[35] <= 32'h03FFF9F8;
                        char22_0[36] <= 32'h01FFF1F8;
                        char22_0[37] <= 32'h003F83F8;
                        char22_0[38] <= 32'h000003F0;
                        char22_0[39] <= 32'h000003F0;
                        char22_0[40] <= 32'h000003F0;
                        char22_0[41] <= 32'h000003F0;
                        char22_0[42] <= 32'h000007E0;
                        char22_0[43] <= 32'h000007E0;
                        char22_0[44] <= 32'h000007C0;
                        char22_0[45] <= 32'h03C007C0;
                        char22_0[46] <= 32'h07C00F80;
                        char22_0[47] <= 32'h0FE00F80;
                        char22_0[48] <= 32'h0FE01F00;
                        char22_0[49] <= 32'h0FE03E00;
                        char22_0[50] <= 32'h07E07E00;
                        char22_0[51] <= 32'h07F1F800;
                        char22_0[52] <= 32'h03FFF000;
                        char22_0[53] <= 32'h00FFC000;
                        char22_0[54] <= 32'h00000000;
                        char22_0[55] <= 32'h00000000;
                        char22_0[56] <= 32'h00000000;
                        char22_0[57] <= 32'h00000000;
                        char22_0[58] <= 32'h00000000;
                        char22_0[59] <= 32'h00000000;
                        char22_0[60] <= 32'h00000000;
                        char22_0[61] <= 32'h00000000;
                        char22_0[62] <= 32'h00000000;
                        char22_0[63] <= 32'h00000000;
                    end//9
                    default: begin
                        char22_0[0] <= char22_0[0];
                        char22_0[1] <= char22_0[1];
                        char22_0[2] <= char22_0[2];
                        char22_0[3] <= char22_0[3];
                        char22_0[4] <= char22_0[4];
                        char22_0[5] <= char22_0[5];
                        char22_0[6] <= char22_0[6];
                        char22_0[7] <= char22_0[7];
                        char22_0[8] <= char22_0[8];
                        char22_0[9] <= char22_0[9];
                        char22_0[10] <= char22_0[10];
                        char22_0[11] <= char22_0[11];
                        char22_0[12] <= char22_0[12];
                        char22_0[13] <= char22_0[13];
                        char22_0[14] <= char22_0[14];
                        char22_0[15] <= char22_0[15];
                        char22_0[16] <= char22_0[16];
                        char22_0[17] <= char22_0[17];
                        char22_0[18] <= char22_0[18];
                        char22_0[19] <= char22_0[19];
                        char22_0[20] <= char22_0[20];
                        char22_0[21] <= char22_0[21];
                        char22_0[22] <= char22_0[22];
                        char22_0[23] <= char22_0[23];
                        char22_0[24] <= char22_0[24];
                        char22_0[25] <= char22_0[25];
                        char22_0[26] <= char22_0[26];
                        char22_0[27] <= char22_0[27];
                        char22_0[28] <= char22_0[28];
                        char22_0[29] <= char22_0[29];
                        char22_0[30] <= char22_0[30];
                        char22_0[31] <= char22_0[31];
                        char22_0[32] <= char22_0[32];
                        char22_0[33] <= char22_0[33];
                        char22_0[34] <= char22_0[34];
                        char22_0[35] <= char22_0[35];
                        char22_0[36] <= char22_0[36];
                        char22_0[37] <= char22_0[37];
                        char22_0[38] <= char22_0[38];
                        char22_0[39] <= char22_0[39];
                        char22_0[40] <= char22_0[40];
                        char22_0[41] <= char22_0[41];
                        char22_0[42] <= char22_0[42];
                        char22_0[43] <= char22_0[43];
                        char22_0[44] <= char22_0[44];
                        char22_0[45] <= char22_0[45];
                        char22_0[46] <= char22_0[46];
                        char22_0[47] <= char22_0[47];
                        char22_0[48] <= char22_0[48];
                        char22_0[49] <= char22_0[49];
                        char22_0[50] <= char22_0[50];
                        char22_0[51] <= char22_0[51];
                        char22_0[52] <= char22_0[52];
                        char22_0[53] <= char22_0[53];
                        char22_0[54] <= char22_0[54];
                        char22_0[55] <= char22_0[55];
                        char22_0[56] <= char22_0[56];
                        char22_0[57] <= char22_0[57];
                        char22_0[58] <= char22_0[58];
                        char22_0[59] <= char22_0[59];
                        char22_0[60] <= char22_0[60];
                        char22_0[61] <= char22_0[61];
                        char22_0[62] <= char22_0[62];
                        char22_0[63] <= char22_0[63];
                    end
                endcase
            
                case((a0 - w1*(a0/w1))/k1)
                        4'd0: begin
                            char22_1[  0] <= 32'h00000000;
                            char22_1[  1] <= 32'h00000000;
                            char22_1[  2] <= 32'h00000000;
                            char22_1[  3] <= 32'h00000000;
                            char22_1[  4] <= 32'h00000000;
                            char22_1[  5] <= 32'h00000000;
                            char22_1[  6] <= 32'h00000000;
                            char22_1[  7] <= 32'h00000000;
                            char22_1[  8] <= 32'h00000000;
                            char22_1[  9] <= 32'h00000000;
                            char22_1[10] <= 32'h000FF000;
                            char22_1[11] <= 32'h003FFC00;
                            char22_1[12] <= 32'h007E7E00;
                            char22_1[13] <= 32'h00F81F00;
                            char22_1[14] <= 32'h01F00F80;
                            char22_1[15] <= 32'h03F00FC0;
                            char22_1[16] <= 32'h03E007C0;
                            char22_1[17] <= 32'h07E007E0;
                            char22_1[18] <= 32'h07C003E0;
                            char22_1[19] <= 32'h0FC003F0;
                            char22_1[20] <= 32'h0FC003F0;
                            char22_1[21] <= 32'h0FC003F0;
                            char22_1[22] <= 32'h1F8001F8;
                            char22_1[23] <= 32'h1F8001F8;
                            char22_1[24] <= 32'h1F8001F8;
                            char22_1[25] <= 32'h1F8001F8;
                            char22_1[26] <= 32'h1F8001F8;
                            char22_1[27] <= 32'h3F8001F8;
                            char22_1[28] <= 32'h3F8001F8;
                            char22_1[29] <= 32'h3F8001F8;
                            char22_1[30] <= 32'h3F8001F8;
                            char22_1[31] <= 32'h3F8001F8;
                            char22_1[32] <= 32'h3F8001F8;
                            char22_1[33] <= 32'h3F8001F8;
                            char22_1[34] <= 32'h3F8001F8;
                            char22_1[35] <= 32'h3F8001F8;
                            char22_1[36] <= 32'h3F8001F8;
                            char22_1[37] <= 32'h1F8001F8;
                            char22_1[38] <= 32'h1F8001F8;
                            char22_1[39] <= 32'h1F8001F8;
                            char22_1[40] <= 32'h1F8001F8;
                            char22_1[41] <= 32'h1F8001F0;
                            char22_1[42] <= 32'h0F8003F0;
                            char22_1[43] <= 32'h0FC003F0;
                            char22_1[44] <= 32'h0FC003F0;
                            char22_1[45] <= 32'h07C003E0;
                            char22_1[46] <= 32'h07E007E0;
                            char22_1[47] <= 32'h03E007C0;
                            char22_1[48] <= 32'h03F00FC0;
                            char22_1[49] <= 32'h01F00F80;
                            char22_1[50] <= 32'h00F81F00;
                            char22_1[51] <= 32'h007E7E00;
                            char22_1[52] <= 32'h003FFC00;
                            char22_1[53] <= 32'h000FF000;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//0
                        4'd1: begin
                            char22_1[  0] <= 32'h00000000;
                            char22_1[  1] <= 32'h00000000;
                            char22_1[  2] <= 32'h00000000;
                            char22_1[  3] <= 32'h00000000;
                            char22_1[  4] <= 32'h00000000;
                            char22_1[  5] <= 32'h00000000;
                            char22_1[  6] <= 32'h00000000;
                            char22_1[  7] <= 32'h00000000;
                            char22_1[  8] <= 32'h00000000;
                            char22_1[  9] <= 32'h00000000;
                            char22_1[10] <= 32'h0000E000;
                            char22_1[11] <= 32'h0001E000;
                            char22_1[12] <= 32'h0003E000;
                            char22_1[13] <= 32'h001FE000;
                            char22_1[14] <= 32'h03FFE000;
                            char22_1[15] <= 32'h03FFE000;
                            char22_1[16] <= 32'h0007E000;
                            char22_1[17] <= 32'h0007E000;
                            char22_1[18] <= 32'h0007E000;
                            char22_1[19] <= 32'h0007E000;
                            char22_1[20] <= 32'h0007E000;
                            char22_1[21] <= 32'h0007E000;
                            char22_1[22] <= 32'h0007E000;
                            char22_1[23] <= 32'h0007E000;
                            char22_1[24] <= 32'h0007E000;
                            char22_1[25] <= 32'h0007E000;
                            char22_1[26] <= 32'h0007E000;
                            char22_1[27] <= 32'h0007E000;
                            char22_1[28] <= 32'h0007E000;
                            char22_1[29] <= 32'h0007E000;
                            char22_1[30] <= 32'h0007E000;
                            char22_1[31] <= 32'h0007E000;
                            char22_1[32] <= 32'h0007E000;
                            char22_1[33] <= 32'h0007E000;
                            char22_1[34] <= 32'h0007E000;
                            char22_1[35] <= 32'h0007E000;
                            char22_1[36] <= 32'h0007E000;
                            char22_1[37] <= 32'h0007E000;
                            char22_1[38] <= 32'h0007E000;
                            char22_1[39] <= 32'h0007E000;
                            char22_1[40] <= 32'h0007E000;
                            char22_1[41] <= 32'h0007E000;
                            char22_1[42] <= 32'h0007E000;
                            char22_1[43] <= 32'h0007E000;
                            char22_1[44] <= 32'h0007E000;
                            char22_1[45] <= 32'h0007E000;
                            char22_1[46] <= 32'h0007E000;
                            char22_1[47] <= 32'h0007E000;
                            char22_1[48] <= 32'h0007E000;
                            char22_1[49] <= 32'h0007E000;
                            char22_1[50] <= 32'h0007E000;
                            char22_1[51] <= 32'h000FF800;
                            char22_1[52] <= 32'h03FFFFC0;
                            char22_1[53] <= 32'h03FFFFC0;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//1
                        4'd2: begin
                            char22_1[  0] <= 32'h00000000;
                            char22_1[  1] <= 32'h00000000;
                            char22_1[  2] <= 32'h00000000;
                            char22_1[  3] <= 32'h00000000;
                            char22_1[  4] <= 32'h00000000;
                            char22_1[  5] <= 32'h00000000;
                            char22_1[  6] <= 32'h00000000;
                            char22_1[  7] <= 32'h00000000;
                            char22_1[  8] <= 32'h00000000;
                            char22_1[  9] <= 32'h00000000;
                            char22_1[10] <= 32'h001FFC00;
                            char22_1[11] <= 32'h007FFF00;
                            char22_1[12] <= 32'h01F83F80;
                            char22_1[13] <= 32'h03E00FC0;
                            char22_1[14] <= 32'h07C007E0;
                            char22_1[15] <= 32'h078007E0;
                            char22_1[16] <= 32'h0F8003F0;
                            char22_1[17] <= 32'h0F8003F0;
                            char22_1[18] <= 32'h1F8003F0;
                            char22_1[19] <= 32'h1F8003F0;
                            char22_1[20] <= 32'h1FC003F0;
                            char22_1[21] <= 32'h1FC003F0;
                            char22_1[22] <= 32'h1FC003F0;
                            char22_1[23] <= 32'h0FC003F0;
                            char22_1[24] <= 32'h07C003F0;
                            char22_1[25] <= 32'h000003E0;
                            char22_1[26] <= 32'h000007E0;
                            char22_1[27] <= 32'h000007E0;
                            char22_1[28] <= 32'h00000FC0;
                            char22_1[29] <= 32'h00000F80;
                            char22_1[30] <= 32'h00001F80;
                            char22_1[31] <= 32'h00003F00;
                            char22_1[32] <= 32'h00003E00;
                            char22_1[33] <= 32'h00007C00;
                            char22_1[34] <= 32'h0000F800;
                            char22_1[35] <= 32'h0001F000;
                            char22_1[36] <= 32'h0003E000;
                            char22_1[37] <= 32'h0007C000;
                            char22_1[38] <= 32'h000F8000;
                            char22_1[39] <= 32'h001F0000;
                            char22_1[40] <= 32'h003E0000;
                            char22_1[41] <= 32'h007C0000;
                            char22_1[42] <= 32'h00F80000;
                            char22_1[43] <= 32'h01F00038;
                            char22_1[44] <= 32'h01E00038;
                            char22_1[45] <= 32'h03C00070;
                            char22_1[46] <= 32'h07800070;
                            char22_1[47] <= 32'h0F8000F0;
                            char22_1[48] <= 32'h0F0000F0;
                            char22_1[49] <= 32'h1E0003F0;
                            char22_1[50] <= 32'h3FFFFFF0;
                            char22_1[51] <= 32'h3FFFFFF0;
                            char22_1[52] <= 32'h3FFFFFE0;
                            char22_1[53] <= 32'h3FFFFFE0;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//2
                        4'd3: begin
                            char22_1[  0] <= 32'h00000000;
                            char22_1[  1] <= 32'h00000000;
                            char22_1[  2] <= 32'h00000000;
                            char22_1[  3] <= 32'h00000000;
                            char22_1[  4] <= 32'h00000000;
                            char22_1[  5] <= 32'h00000000;
                            char22_1[  6] <= 32'h00000000;
                            char22_1[  7] <= 32'h00000000;
                            char22_1[  8] <= 32'h00000000;
                            char22_1[  9] <= 32'h00000000;
                            char22_1[10] <= 32'h003FF000;
                            char22_1[11] <= 32'h00FFFC00;
                            char22_1[12] <= 32'h01F07E00;
                            char22_1[13] <= 32'h03C03F00;
                            char22_1[14] <= 32'h07801F80;
                            char22_1[15] <= 32'h0F800FC0;
                            char22_1[16] <= 32'h0F800FC0;
                            char22_1[17] <= 32'h0F8007E0;
                            char22_1[18] <= 32'h0FC007E0;
                            char22_1[19] <= 32'h0FC007E0;
                            char22_1[20] <= 32'h0FC007E0;
                            char22_1[21] <= 32'h07C007E0;
                            char22_1[22] <= 32'h000007E0;
                            char22_1[23] <= 32'h000007E0;
                            char22_1[24] <= 32'h000007C0;
                            char22_1[25] <= 32'h00000FC0;
                            char22_1[26] <= 32'h00000F80;
                            char22_1[27] <= 32'h00001F00;
                            char22_1[28] <= 32'h00007E00;
                            char22_1[29] <= 32'h0003FC00;
                            char22_1[30] <= 32'h001FF000;
                            char22_1[31] <= 32'h001FFC00;
                            char22_1[32] <= 32'h0000FF00;
                            char22_1[33] <= 32'h00001F80;
                            char22_1[34] <= 32'h00000FC0;
                            char22_1[35] <= 32'h000007E0;
                            char22_1[36] <= 32'h000003E0;
                            char22_1[37] <= 32'h000003F0;
                            char22_1[38] <= 32'h000003F0;
                            char22_1[39] <= 32'h000001F0;
                            char22_1[40] <= 32'h000001F8;
                            char22_1[41] <= 32'h000001F8;
                            char22_1[42] <= 32'h078001F8;
                            char22_1[43] <= 32'h0FC001F8;
                            char22_1[44] <= 32'h1FC001F8;
                            char22_1[45] <= 32'h1FC003F0;
                            char22_1[46] <= 32'h1FC003F0;
                            char22_1[47] <= 32'h1FC003E0;
                            char22_1[48] <= 32'h0F8007E0;
                            char22_1[49] <= 32'h0F8007C0;
                            char22_1[50] <= 32'h07C01F80;
                            char22_1[51] <= 32'h03F07F00;
                            char22_1[52] <= 32'h01FFFE00;
                            char22_1[53] <= 32'h003FF000;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//3
                        4'd4: begin
                            char22_1[  0] <= 32'h00000000;
                            char22_1[  1] <= 32'h00000000;
                            char22_1[  2] <= 32'h00000000;
                            char22_1[  3] <= 32'h00000000;
                            char22_1[  4] <= 32'h00000000;
                            char22_1[  5] <= 32'h00000000;
                            char22_1[  6] <= 32'h00000000;
                            char22_1[  7] <= 32'h00000000;
                            char22_1[  8] <= 32'h00000000;
                            char22_1[  9] <= 32'h00000000;
                            char22_1[10] <= 32'h00001F00;
                            char22_1[11] <= 32'h00001F00;
                            char22_1[12] <= 32'h00003F00;
                            char22_1[13] <= 32'h00003F00;
                            char22_1[14] <= 32'h00007F00;
                            char22_1[15] <= 32'h0000FF00;
                            char22_1[16] <= 32'h0000FF00;
                            char22_1[17] <= 32'h0001FF00;
                            char22_1[18] <= 32'h0003FF00;
                            char22_1[19] <= 32'h0003BF00;
                            char22_1[20] <= 32'h0007BF00;
                            char22_1[21] <= 32'h00073F00;
                            char22_1[22] <= 32'h000F3F00;
                            char22_1[23] <= 32'h001E3F00;
                            char22_1[24] <= 32'h001C3F00;
                            char22_1[25] <= 32'h003C3F00;
                            char22_1[26] <= 32'h00783F00;
                            char22_1[27] <= 32'h00783F00;
                            char22_1[28] <= 32'h00F03F00;
                            char22_1[29] <= 32'h00E03F00;
                            char22_1[30] <= 32'h01E03F00;
                            char22_1[31] <= 32'h03C03F00;
                            char22_1[32] <= 32'h03803F00;
                            char22_1[33] <= 32'h07803F00;
                            char22_1[34] <= 32'h0F003F00;
                            char22_1[35] <= 32'h0F003F00;
                            char22_1[36] <= 32'h1E003F00;
                            char22_1[37] <= 32'h1C003F00;
                            char22_1[38] <= 32'h3C003F00;
                            char22_1[39] <= 32'h7FFFFFFE;
                            char22_1[40] <= 32'h7FFFFFFE;
                            char22_1[41] <= 32'h00003F00;
                            char22_1[42] <= 32'h00003F00;
                            char22_1[43] <= 32'h00003F00;
                            char22_1[44] <= 32'h00003F00;
                            char22_1[45] <= 32'h00003F00;
                            char22_1[46] <= 32'h00003F00;
                            char22_1[47] <= 32'h00003F00;
                            char22_1[48] <= 32'h00003F00;
                            char22_1[49] <= 32'h00003F00;
                            char22_1[50] <= 32'h00003F00;
                            char22_1[51] <= 32'h00007F80;
                            char22_1[52] <= 32'h000FFFFC;
                            char22_1[53] <= 32'h000FFFFC;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//4
                        4'd5: begin
                            char22_1[  0] <= 32'h00000000;
                            char22_1[  1] <= 32'h00000000;
                            char22_1[  2] <= 32'h00000000;
                            char22_1[  3] <= 32'h00000000;
                            char22_1[  4] <= 32'h00000000;
                            char22_1[  5] <= 32'h00000000;
                            char22_1[  6] <= 32'h00000000;
                            char22_1[  7] <= 32'h00000000;
                            char22_1[  8] <= 32'h00000000;
                            char22_1[  9] <= 32'h00000000;
                            char22_1[10] <= 32'h00000000;
                            char22_1[11] <= 32'h03FFFFF0;
                            char22_1[12] <= 32'h03FFFFF0;
                            char22_1[13] <= 32'h03FFFFF0;
                            char22_1[14] <= 32'h03FFFFE0;
                            char22_1[15] <= 32'h03800000;
                            char22_1[16] <= 32'h03800000;
                            char22_1[17] <= 32'h03800000;
                            char22_1[18] <= 32'h03800000;
                            char22_1[19] <= 32'h03800000;
                            char22_1[20] <= 32'h07800000;
                            char22_1[21] <= 32'h07800000;
                            char22_1[22] <= 32'h07800000;
                            char22_1[23] <= 32'h07800000;
                            char22_1[24] <= 32'h07800000;
                            char22_1[25] <= 32'h07800000;
                            char22_1[26] <= 32'h078FF800;
                            char22_1[27] <= 32'h073FFE00;
                            char22_1[28] <= 32'h077FFF80;
                            char22_1[29] <= 32'h07FC3F80;
                            char22_1[30] <= 32'h07E00FC0;
                            char22_1[31] <= 32'h07C007E0;
                            char22_1[32] <= 32'h078007E0;
                            char22_1[33] <= 32'h078003F0;
                            char22_1[34] <= 32'h000003F0;
                            char22_1[35] <= 32'h000001F0;
                            char22_1[36] <= 32'h000001F8;
                            char22_1[37] <= 32'h000001F8;
                            char22_1[38] <= 32'h000001F8;
                            char22_1[39] <= 32'h000001F8;
                            char22_1[40] <= 32'h000001F8;
                            char22_1[41] <= 32'h078001F8;
                            char22_1[42] <= 32'h0FC001F8;
                            char22_1[43] <= 32'h1FC001F0;
                            char22_1[44] <= 32'h1FC001F0;
                            char22_1[45] <= 32'h1FC003F0;
                            char22_1[46] <= 32'h1F8003F0;
                            char22_1[47] <= 32'h1F8003E0;
                            char22_1[48] <= 32'h0F8007E0;
                            char22_1[49] <= 32'h078007C0;
                            char22_1[50] <= 32'h07C01F80;
                            char22_1[51] <= 32'h03F83F00;
                            char22_1[52] <= 32'h00FFFE00;
                            char22_1[53] <= 32'h003FF800;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//5
                        4'd6: begin
                            char22_1[0] <= 32'h00000000;
                            char22_1[1] <= 32'h00000000;
                            char22_1[2] <= 32'h00000000;
                            char22_1[3] <= 32'h00000000;
                            char22_1[4] <= 32'h00000000;
                            char22_1[5] <= 32'h00000000;
                            char22_1[6] <= 32'h00000000;
                            char22_1[7] <= 32'h00000000;
                            char22_1[8] <= 32'h00000000;
                            char22_1[9] <= 32'h00000000;
                            char22_1[10] <= 32'h0007FE00;
                            char22_1[11] <= 32'h001FFF80;
                            char22_1[12] <= 32'h003F0FC0;
                            char22_1[13] <= 32'h007C07C0;
                            char22_1[14] <= 32'h00F807E0;
                            char22_1[15] <= 32'h01F007E0;
                            char22_1[16] <= 32'h03E007E0;
                            char22_1[17] <= 32'h03C007E0;
                            char22_1[18] <= 32'h07C003C0;
                            char22_1[19] <= 32'h07C00000;
                            char22_1[20] <= 32'h0FC00000;
                            char22_1[21] <= 32'h0F800000;
                            char22_1[22] <= 32'h0F800000;
                            char22_1[23] <= 32'h1F800000;
                            char22_1[24] <= 32'h1F800000;
                            char22_1[25] <= 32'h1F800000;
                            char22_1[26] <= 32'h1F87FE00;
                            char22_1[27] <= 32'h1F9FFF80;
                            char22_1[28] <= 32'h1FBFFFC0;
                            char22_1[29] <= 32'h3FFE1FC0;
                            char22_1[30] <= 32'h3FF807E0;
                            char22_1[31] <= 32'h3FE003F0;
                            char22_1[32] <= 32'h3FE003F0;
                            char22_1[33] <= 32'h3FC001F8;
                            char22_1[34] <= 32'h3F8001F8;
                            char22_1[35] <= 32'h3F8001F8;
                            char22_1[36] <= 32'h3F8000F8;
                            char22_1[37] <= 32'h3F8000F8;
                            char22_1[38] <= 32'h3F8000F8;
                            char22_1[39] <= 32'h1F8000F8;
                            char22_1[40] <= 32'h1F8000F8;
                            char22_1[41] <= 32'h1F8000F8;
                            char22_1[42] <= 32'h1F8000F8;
                            char22_1[43] <= 32'h1F8000F8;
                            char22_1[44] <= 32'h0FC001F8;
                            char22_1[45] <= 32'h0FC001F8;
                            char22_1[46] <= 32'h0FC001F0;
                            char22_1[47] <= 32'h07E001F0;
                            char22_1[48] <= 32'h03E003E0;
                            char22_1[49] <= 32'h03F003E0;
                            char22_1[50] <= 32'h01F807C0;
                            char22_1[51] <= 32'h00FE1F80;
                            char22_1[52] <= 32'h007FFE00;
                            char22_1[53] <= 32'h001FF800;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//6
                        4'd7: begin
                            char22_1[0] <= 32'h00000000;
                            char22_1[1] <= 32'h00000000;
                            char22_1[2] <= 32'h00000000;
                            char22_1[3] <= 32'h00000000;
                            char22_1[4] <= 32'h00000000;
                            char22_1[5] <= 32'h00000000;
                            char22_1[6] <= 32'h00000000;
                            char22_1[7] <= 32'h00000000;
                            char22_1[8] <= 32'h00000000;
                            char22_1[9] <= 32'h00000000;
                            char22_1[10] <= 32'h00000000;
                            char22_1[11] <= 32'h07FFFFF8;
                            char22_1[12] <= 32'h07FFFFF8;
                            char22_1[13] <= 32'h07FFFFF8;
                            char22_1[14] <= 32'h0FFFFFF0;
                            char22_1[15] <= 32'h0FC000E0;
                            char22_1[16] <= 32'h0F8001E0;
                            char22_1[17] <= 32'h0F0001C0;
                            char22_1[18] <= 32'h0E0003C0;
                            char22_1[19] <= 32'h0E000780;
                            char22_1[20] <= 32'h1E000780;
                            char22_1[21] <= 32'h1C000F00;
                            char22_1[22] <= 32'h00000F00;
                            char22_1[23] <= 32'h00001E00;
                            char22_1[24] <= 32'h00001E00;
                            char22_1[25] <= 32'h00003C00;
                            char22_1[26] <= 32'h00003C00;
                            char22_1[27] <= 32'h00007800;
                            char22_1[28] <= 32'h00007800;
                            char22_1[29] <= 32'h0000F800;
                            char22_1[30] <= 32'h0000F000;
                            char22_1[31] <= 32'h0001F000;
                            char22_1[32] <= 32'h0001E000;
                            char22_1[33] <= 32'h0003E000;
                            char22_1[34] <= 32'h0003E000;
                            char22_1[35] <= 32'h0003E000;
                            char22_1[36] <= 32'h0007C000;
                            char22_1[37] <= 32'h0007C000;
                            char22_1[38] <= 32'h0007C000;
                            char22_1[39] <= 32'h000FC000;
                            char22_1[40] <= 32'h000FC000;
                            char22_1[41] <= 32'h000FC000;
                            char22_1[42] <= 32'h000FC000;
                            char22_1[43] <= 32'h001FC000;
                            char22_1[44] <= 32'h001FC000;
                            char22_1[45] <= 32'h001FC000;
                            char22_1[46] <= 32'h001FC000;
                            char22_1[47] <= 32'h001FC000;
                            char22_1[48] <= 32'h001FC000;
                            char22_1[49] <= 32'h001FC000;
                            char22_1[50] <= 32'h001FC000;
                            char22_1[51] <= 32'h001FC000;
                            char22_1[52] <= 32'h001FC000;
                            char22_1[53] <= 32'h000F8000;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//7
                        4'd8: begin
                            char22_1[0] <= 32'h00000000;
                            char22_1[1] <= 32'h00000000;
                            char22_1[2] <= 32'h00000000;
                            char22_1[3] <= 32'h00000000;
                            char22_1[4] <= 32'h00000000;
                            char22_1[5] <= 32'h00000000;
                            char22_1[6] <= 32'h00000000;
                            char22_1[7] <= 32'h00000000;
                            char22_1[8] <= 32'h00000000;
                            char22_1[9] <= 32'h00000000;
                            char22_1[10] <= 32'h003FF800;
                            char22_1[11] <= 32'h00FFFE00;
                            char22_1[12] <= 32'h01F81F80;
                            char22_1[13] <= 32'h03E00FC0;
                            char22_1[14] <= 32'h07C003E0;
                            char22_1[15] <= 32'h0F8003E0;
                            char22_1[16] <= 32'h0F8001F0;
                            char22_1[17] <= 32'h1F0001F0;
                            char22_1[18] <= 32'h1F0001F0;
                            char22_1[19] <= 32'h1F0001F0;
                            char22_1[20] <= 32'h1F0001F0;
                            char22_1[21] <= 32'h1F0001F0;
                            char22_1[22] <= 32'h1F8001F0;
                            char22_1[23] <= 32'h1FC001F0;
                            char22_1[24] <= 32'h0FC001F0;
                            char22_1[25] <= 32'h0FF003E0;
                            char22_1[26] <= 32'h07F803C0;
                            char22_1[27] <= 32'h03FE0F80;
                            char22_1[28] <= 32'h01FF9F00;
                            char22_1[29] <= 32'h00FFFE00;
                            char22_1[30] <= 32'h003FF800;
                            char22_1[31] <= 32'h007FFC00;
                            char22_1[32] <= 32'h01F7FF00;
                            char22_1[33] <= 32'h03E1FF80;
                            char22_1[34] <= 32'h07C07FC0;
                            char22_1[35] <= 32'h0F801FE0;
                            char22_1[36] <= 32'h0F800FE0;
                            char22_1[37] <= 32'h1F0007F0;
                            char22_1[38] <= 32'h1F0003F0;
                            char22_1[39] <= 32'h3E0001F8;
                            char22_1[40] <= 32'h3E0001F8;
                            char22_1[41] <= 32'h3E0001F8;
                            char22_1[42] <= 32'h3E0000F8;
                            char22_1[43] <= 32'h3E0000F8;
                            char22_1[44] <= 32'h3E0000F8;
                            char22_1[45] <= 32'h3E0000F8;
                            char22_1[46] <= 32'h1F0001F0;
                            char22_1[47] <= 32'h1F0001F0;
                            char22_1[48] <= 32'h0F8003E0;
                            char22_1[49] <= 32'h0FC003E0;
                            char22_1[50] <= 32'h07E007C0;
                            char22_1[51] <= 32'h01F83F80;
                            char22_1[52] <= 32'h00FFFE00;
                            char22_1[53] <= 32'h003FF800;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//8
                        4'd9: begin
                            char22_1[0] <= 32'h00000000;
                            char22_1[1] <= 32'h00000000;
                            char22_1[2] <= 32'h00000000;
                            char22_1[3] <= 32'h00000000;
                            char22_1[4] <= 32'h00000000;
                            char22_1[5] <= 32'h00000000;
                            char22_1[6] <= 32'h00000000;
                            char22_1[7] <= 32'h00000000;
                            char22_1[8] <= 32'h00000000;
                            char22_1[9] <= 32'h00000000;
                            char22_1[10] <= 32'h003FF000;
                            char22_1[11] <= 32'h00FFFC00;
                            char22_1[12] <= 32'h01F83F00;
                            char22_1[13] <= 32'h03E01F80;
                            char22_1[14] <= 32'h07C00F80;
                            char22_1[15] <= 32'h0FC007C0;
                            char22_1[16] <= 32'h0F8003E0;
                            char22_1[17] <= 32'h1F8003E0;
                            char22_1[18] <= 32'h1F0003F0;
                            char22_1[19] <= 32'h1F0003F0;
                            char22_1[20] <= 32'h3F0001F0;
                            char22_1[21] <= 32'h3F0001F0;
                            char22_1[22] <= 32'h3F0001F8;
                            char22_1[23] <= 32'h3F0001F8;
                            char22_1[24] <= 32'h3F0001F8;
                            char22_1[25] <= 32'h3F0001F8;
                            char22_1[26] <= 32'h3F0001F8;
                            char22_1[27] <= 32'h3F0001F8;
                            char22_1[28] <= 32'h3F0003F8;
                            char22_1[29] <= 32'h1F8003F8;
                            char22_1[30] <= 32'h1F8007F8;
                            char22_1[31] <= 32'h1F800FF8;
                            char22_1[32] <= 32'h0FC01FF8;
                            char22_1[33] <= 32'h0FE03FF8;
                            char22_1[34] <= 32'h07F8FDF8;
                            char22_1[35] <= 32'h03FFF9F8;
                            char22_1[36] <= 32'h01FFF1F8;
                            char22_1[37] <= 32'h003F83F8;
                            char22_1[38] <= 32'h000003F0;
                            char22_1[39] <= 32'h000003F0;
                            char22_1[40] <= 32'h000003F0;
                            char22_1[41] <= 32'h000003F0;
                            char22_1[42] <= 32'h000007E0;
                            char22_1[43] <= 32'h000007E0;
                            char22_1[44] <= 32'h000007C0;
                            char22_1[45] <= 32'h03C007C0;
                            char22_1[46] <= 32'h07C00F80;
                            char22_1[47] <= 32'h0FE00F80;
                            char22_1[48] <= 32'h0FE01F00;
                            char22_1[49] <= 32'h0FE03E00;
                            char22_1[50] <= 32'h07E07E00;
                            char22_1[51] <= 32'h07F1F800;
                            char22_1[52] <= 32'h03FFF000;
                            char22_1[53] <= 32'h00FFC000;
                            char22_1[54] <= 32'h00000000;
                            char22_1[55] <= 32'h00000000;
                            char22_1[56] <= 32'h00000000;
                            char22_1[57] <= 32'h00000000;
                            char22_1[58] <= 32'h00000000;
                            char22_1[59] <= 32'h00000000;
                            char22_1[60] <= 32'h00000000;
                            char22_1[61] <= 32'h00000000;
                            char22_1[62] <= 32'h00000000;
                            char22_1[63] <= 32'h00000000;
                        end//9
                        default: begin
                            char22_1[0] <= char22_1[0];
                            char22_1[1] <= char22_1[1];
                            char22_1[2] <= char22_1[2];
                            char22_1[3] <= char22_1[3];
                            char22_1[4] <= char22_1[4];
                            char22_1[5] <= char22_1[5];
                            char22_1[6] <= char22_1[6];
                            char22_1[7] <= char22_1[7];
                            char22_1[8] <= char22_1[8];
                            char22_1[9] <= char22_1[9];
                            char22_1[10] <= char22_1[10];
                            char22_1[11] <= char22_1[11];
                            char22_1[12] <= char22_1[12];
                            char22_1[13] <= char22_1[13];
                            char22_1[14] <= char22_1[14];
                            char22_1[15] <= char22_1[15];
                            char22_1[16] <= char22_1[16];
                            char22_1[17] <= char22_1[17];
                            char22_1[18] <= char22_1[18];
                            char22_1[19] <= char22_1[19];
                            char22_1[20] <= char22_1[20];
                            char22_1[21] <= char22_1[21];
                            char22_1[22] <= char22_1[22];
                            char22_1[23] <= char22_1[23];
                            char22_1[24] <= char22_1[24];
                            char22_1[25] <= char22_1[25];
                            char22_1[26] <= char22_1[26];
                            char22_1[27] <= char22_1[27];
                            char22_1[28] <= char22_1[28];
                            char22_1[29] <= char22_1[29];
                            char22_1[30] <= char22_1[30];
                            char22_1[31] <= char22_1[31];
                            char22_1[32] <= char22_1[32];
                            char22_1[33] <= char22_1[33];
                            char22_1[34] <= char22_1[34];
                            char22_1[35] <= char22_1[35];
                            char22_1[36] <= char22_1[36];
                            char22_1[37] <= char22_1[37];
                            char22_1[38] <= char22_1[38];
                            char22_1[39] <= char22_1[39];
                            char22_1[40] <= char22_1[40];
                            char22_1[41] <= char22_1[41];
                            char22_1[42] <= char22_1[42];
                            char22_1[43] <= char22_1[43];
                            char22_1[44] <= char22_1[44];
                            char22_1[45] <= char22_1[45];
                            char22_1[46] <= char22_1[46];
                            char22_1[47] <= char22_1[47];
                            char22_1[48] <= char22_1[48];
                            char22_1[49] <= char22_1[49];
                            char22_1[50] <= char22_1[50];
                            char22_1[51] <= char22_1[51];
                            char22_1[52] <= char22_1[52];
                            char22_1[53] <= char22_1[53];
                            char22_1[54] <= char22_1[54];
                            char22_1[55] <= char22_1[55];
                            char22_1[56] <= char22_1[56];
                            char22_1[57] <= char22_1[57];
                            char22_1[58] <= char22_1[58];
                            char22_1[59] <= char22_1[59];
                            char22_1[60] <= char22_1[60];
                            char22_1[61] <= char22_1[61];
                            char22_1[62] <= char22_1[62];
                            char22_1[63] <= char22_1[63];
                        end
                    endcase
            
                case((a0 - k1*(a0/k1))/h1)
                            4'd0: begin
                                char22_2[  0] <= 32'h00000000;
                                char22_2[  1] <= 32'h00000000;
                                char22_2[  2] <= 32'h00000000;
                                char22_2[  3] <= 32'h00000000;
                                char22_2[  4] <= 32'h00000000;
                                char22_2[  5] <= 32'h00000000;
                                char22_2[  6] <= 32'h00000000;
                                char22_2[  7] <= 32'h00000000;
                                char22_2[  8] <= 32'h00000000;
                                char22_2[  9] <= 32'h00000000;
                                char22_2[10] <= 32'h000FF000;
                                char22_2[11] <= 32'h003FFC00;
                                char22_2[12] <= 32'h007E7E00;
                                char22_2[13] <= 32'h00F81F00;
                                char22_2[14] <= 32'h01F00F80;
                                char22_2[15] <= 32'h03F00FC0;
                                char22_2[16] <= 32'h03E007C0;
                                char22_2[17] <= 32'h07E007E0;
                                char22_2[18] <= 32'h07C003E0;
                                char22_2[19] <= 32'h0FC003F0;
                                char22_2[20] <= 32'h0FC003F0;
                                char22_2[21] <= 32'h0FC003F0;
                                char22_2[22] <= 32'h1F8001F8;
                                char22_2[23] <= 32'h1F8001F8;
                                char22_2[24] <= 32'h1F8001F8;
                                char22_2[25] <= 32'h1F8001F8;
                                char22_2[26] <= 32'h1F8001F8;
                                char22_2[27] <= 32'h3F8001F8;
                                char22_2[28] <= 32'h3F8001F8;
                                char22_2[29] <= 32'h3F8001F8;
                                char22_2[30] <= 32'h3F8001F8;
                                char22_2[31] <= 32'h3F8001F8;
                                char22_2[32] <= 32'h3F8001F8;
                                char22_2[33] <= 32'h3F8001F8;
                                char22_2[34] <= 32'h3F8001F8;
                                char22_2[35] <= 32'h3F8001F8;
                                char22_2[36] <= 32'h3F8001F8;
                                char22_2[37] <= 32'h1F8001F8;
                                char22_2[38] <= 32'h1F8001F8;
                                char22_2[39] <= 32'h1F8001F8;
                                char22_2[40] <= 32'h1F8001F8;
                                char22_2[41] <= 32'h1F8001F0;
                                char22_2[42] <= 32'h0F8003F0;
                                char22_2[43] <= 32'h0FC003F0;
                                char22_2[44] <= 32'h0FC003F0;
                                char22_2[45] <= 32'h07C003E0;
                                char22_2[46] <= 32'h07E007E0;
                                char22_2[47] <= 32'h03E007C0;
                                char22_2[48] <= 32'h03F00FC0;
                                char22_2[49] <= 32'h01F00F80;
                                char22_2[50] <= 32'h00F81F00;
                                char22_2[51] <= 32'h007E7E00;
                                char22_2[52] <= 32'h003FFC00;
                                char22_2[53] <= 32'h000FF000;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//0
                            4'd1: begin
                                char22_2[  0] <= 32'h00000000;
                                char22_2[  1] <= 32'h00000000;
                                char22_2[  2] <= 32'h00000000;
                                char22_2[  3] <= 32'h00000000;
                                char22_2[  4] <= 32'h00000000;
                                char22_2[  5] <= 32'h00000000;
                                char22_2[  6] <= 32'h00000000;
                                char22_2[  7] <= 32'h00000000;
                                char22_2[  8] <= 32'h00000000;
                                char22_2[  9] <= 32'h00000000;
                                char22_2[10] <= 32'h0000E000;
                                char22_2[11] <= 32'h0001E000;
                                char22_2[12] <= 32'h0003E000;
                                char22_2[13] <= 32'h001FE000;
                                char22_2[14] <= 32'h03FFE000;
                                char22_2[15] <= 32'h03FFE000;
                                char22_2[16] <= 32'h0007E000;
                                char22_2[17] <= 32'h0007E000;
                                char22_2[18] <= 32'h0007E000;
                                char22_2[19] <= 32'h0007E000;
                                char22_2[20] <= 32'h0007E000;
                                char22_2[21] <= 32'h0007E000;
                                char22_2[22] <= 32'h0007E000;
                                char22_2[23] <= 32'h0007E000;
                                char22_2[24] <= 32'h0007E000;
                                char22_2[25] <= 32'h0007E000;
                                char22_2[26] <= 32'h0007E000;
                                char22_2[27] <= 32'h0007E000;
                                char22_2[28] <= 32'h0007E000;
                                char22_2[29] <= 32'h0007E000;
                                char22_2[30] <= 32'h0007E000;
                                char22_2[31] <= 32'h0007E000;
                                char22_2[32] <= 32'h0007E000;
                                char22_2[33] <= 32'h0007E000;
                                char22_2[34] <= 32'h0007E000;
                                char22_2[35] <= 32'h0007E000;
                                char22_2[36] <= 32'h0007E000;
                                char22_2[37] <= 32'h0007E000;
                                char22_2[38] <= 32'h0007E000;
                                char22_2[39] <= 32'h0007E000;
                                char22_2[40] <= 32'h0007E000;
                                char22_2[41] <= 32'h0007E000;
                                char22_2[42] <= 32'h0007E000;
                                char22_2[43] <= 32'h0007E000;
                                char22_2[44] <= 32'h0007E000;
                                char22_2[45] <= 32'h0007E000;
                                char22_2[46] <= 32'h0007E000;
                                char22_2[47] <= 32'h0007E000;
                                char22_2[48] <= 32'h0007E000;
                                char22_2[49] <= 32'h0007E000;
                                char22_2[50] <= 32'h0007E000;
                                char22_2[51] <= 32'h000FF800;
                                char22_2[52] <= 32'h03FFFFC0;
                                char22_2[53] <= 32'h03FFFFC0;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//1
                            4'd2: begin
                                char22_2[  0] <= 32'h00000000;
                                char22_2[  1] <= 32'h00000000;
                                char22_2[  2] <= 32'h00000000;
                                char22_2[  3] <= 32'h00000000;
                                char22_2[  4] <= 32'h00000000;
                                char22_2[  5] <= 32'h00000000;
                                char22_2[  6] <= 32'h00000000;
                                char22_2[  7] <= 32'h00000000;
                                char22_2[  8] <= 32'h00000000;
                                char22_2[  9] <= 32'h00000000;
                                char22_2[10] <= 32'h001FFC00;
                                char22_2[11] <= 32'h007FFF00;
                                char22_2[12] <= 32'h01F83F80;
                                char22_2[13] <= 32'h03E00FC0;
                                char22_2[14] <= 32'h07C007E0;
                                char22_2[15] <= 32'h078007E0;
                                char22_2[16] <= 32'h0F8003F0;
                                char22_2[17] <= 32'h0F8003F0;
                                char22_2[18] <= 32'h1F8003F0;
                                char22_2[19] <= 32'h1F8003F0;
                                char22_2[20] <= 32'h1FC003F0;
                                char22_2[21] <= 32'h1FC003F0;
                                char22_2[22] <= 32'h1FC003F0;
                                char22_2[23] <= 32'h0FC003F0;
                                char22_2[24] <= 32'h07C003F0;
                                char22_2[25] <= 32'h000003E0;
                                char22_2[26] <= 32'h000007E0;
                                char22_2[27] <= 32'h000007E0;
                                char22_2[28] <= 32'h00000FC0;
                                char22_2[29] <= 32'h00000F80;
                                char22_2[30] <= 32'h00001F80;
                                char22_2[31] <= 32'h00003F00;
                                char22_2[32] <= 32'h00003E00;
                                char22_2[33] <= 32'h00007C00;
                                char22_2[34] <= 32'h0000F800;
                                char22_2[35] <= 32'h0001F000;
                                char22_2[36] <= 32'h0003E000;
                                char22_2[37] <= 32'h0007C000;
                                char22_2[38] <= 32'h000F8000;
                                char22_2[39] <= 32'h001F0000;
                                char22_2[40] <= 32'h003E0000;
                                char22_2[41] <= 32'h007C0000;
                                char22_2[42] <= 32'h00F80000;
                                char22_2[43] <= 32'h01F00038;
                                char22_2[44] <= 32'h01E00038;
                                char22_2[45] <= 32'h03C00070;
                                char22_2[46] <= 32'h07800070;
                                char22_2[47] <= 32'h0F8000F0;
                                char22_2[48] <= 32'h0F0000F0;
                                char22_2[49] <= 32'h1E0003F0;
                                char22_2[50] <= 32'h3FFFFFF0;
                                char22_2[51] <= 32'h3FFFFFF0;
                                char22_2[52] <= 32'h3FFFFFE0;
                                char22_2[53] <= 32'h3FFFFFE0;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//2
                            4'd3: begin
                                char22_2[  0] <= 32'h00000000;
                                char22_2[  1] <= 32'h00000000;
                                char22_2[  2] <= 32'h00000000;
                                char22_2[  3] <= 32'h00000000;
                                char22_2[  4] <= 32'h00000000;
                                char22_2[  5] <= 32'h00000000;
                                char22_2[  6] <= 32'h00000000;
                                char22_2[  7] <= 32'h00000000;
                                char22_2[  8] <= 32'h00000000;
                                char22_2[  9] <= 32'h00000000;
                                char22_2[10] <= 32'h003FF000;
                                char22_2[11] <= 32'h00FFFC00;
                                char22_2[12] <= 32'h01F07E00;
                                char22_2[13] <= 32'h03C03F00;
                                char22_2[14] <= 32'h07801F80;
                                char22_2[15] <= 32'h0F800FC0;
                                char22_2[16] <= 32'h0F800FC0;
                                char22_2[17] <= 32'h0F8007E0;
                                char22_2[18] <= 32'h0FC007E0;
                                char22_2[19] <= 32'h0FC007E0;
                                char22_2[20] <= 32'h0FC007E0;
                                char22_2[21] <= 32'h07C007E0;
                                char22_2[22] <= 32'h000007E0;
                                char22_2[23] <= 32'h000007E0;
                                char22_2[24] <= 32'h000007C0;
                                char22_2[25] <= 32'h00000FC0;
                                char22_2[26] <= 32'h00000F80;
                                char22_2[27] <= 32'h00001F00;
                                char22_2[28] <= 32'h00007E00;
                                char22_2[29] <= 32'h0003FC00;
                                char22_2[30] <= 32'h001FF000;
                                char22_2[31] <= 32'h001FFC00;
                                char22_2[32] <= 32'h0000FF00;
                                char22_2[33] <= 32'h00001F80;
                                char22_2[34] <= 32'h00000FC0;
                                char22_2[35] <= 32'h000007E0;
                                char22_2[36] <= 32'h000003E0;
                                char22_2[37] <= 32'h000003F0;
                                char22_2[38] <= 32'h000003F0;
                                char22_2[39] <= 32'h000001F0;
                                char22_2[40] <= 32'h000001F8;
                                char22_2[41] <= 32'h000001F8;
                                char22_2[42] <= 32'h078001F8;
                                char22_2[43] <= 32'h0FC001F8;
                                char22_2[44] <= 32'h1FC001F8;
                                char22_2[45] <= 32'h1FC003F0;
                                char22_2[46] <= 32'h1FC003F0;
                                char22_2[47] <= 32'h1FC003E0;
                                char22_2[48] <= 32'h0F8007E0;
                                char22_2[49] <= 32'h0F8007C0;
                                char22_2[50] <= 32'h07C01F80;
                                char22_2[51] <= 32'h03F07F00;
                                char22_2[52] <= 32'h01FFFE00;
                                char22_2[53] <= 32'h003FF000;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//3
                            4'd4: begin
                                char22_2[  0] <= 32'h00000000;
                                char22_2[  1] <= 32'h00000000;
                                char22_2[  2] <= 32'h00000000;
                                char22_2[  3] <= 32'h00000000;
                                char22_2[  4] <= 32'h00000000;
                                char22_2[  5] <= 32'h00000000;
                                char22_2[  6] <= 32'h00000000;
                                char22_2[  7] <= 32'h00000000;
                                char22_2[  8] <= 32'h00000000;
                                char22_2[  9] <= 32'h00000000;
                                char22_2[10] <= 32'h00001F00;
                                char22_2[11] <= 32'h00001F00;
                                char22_2[12] <= 32'h00003F00;
                                char22_2[13] <= 32'h00003F00;
                                char22_2[14] <= 32'h00007F00;
                                char22_2[15] <= 32'h0000FF00;
                                char22_2[16] <= 32'h0000FF00;
                                char22_2[17] <= 32'h0001FF00;
                                char22_2[18] <= 32'h0003FF00;
                                char22_2[19] <= 32'h0003BF00;
                                char22_2[20] <= 32'h0007BF00;
                                char22_2[21] <= 32'h00073F00;
                                char22_2[22] <= 32'h000F3F00;
                                char22_2[23] <= 32'h001E3F00;
                                char22_2[24] <= 32'h001C3F00;
                                char22_2[25] <= 32'h003C3F00;
                                char22_2[26] <= 32'h00783F00;
                                char22_2[27] <= 32'h00783F00;
                                char22_2[28] <= 32'h00F03F00;
                                char22_2[29] <= 32'h00E03F00;
                                char22_2[30] <= 32'h01E03F00;
                                char22_2[31] <= 32'h03C03F00;
                                char22_2[32] <= 32'h03803F00;
                                char22_2[33] <= 32'h07803F00;
                                char22_2[34] <= 32'h0F003F00;
                                char22_2[35] <= 32'h0F003F00;
                                char22_2[36] <= 32'h1E003F00;
                                char22_2[37] <= 32'h1C003F00;
                                char22_2[38] <= 32'h3C003F00;
                                char22_2[39] <= 32'h7FFFFFFE;
                                char22_2[40] <= 32'h7FFFFFFE;
                                char22_2[41] <= 32'h00003F00;
                                char22_2[42] <= 32'h00003F00;
                                char22_2[43] <= 32'h00003F00;
                                char22_2[44] <= 32'h00003F00;
                                char22_2[45] <= 32'h00003F00;
                                char22_2[46] <= 32'h00003F00;
                                char22_2[47] <= 32'h00003F00;
                                char22_2[48] <= 32'h00003F00;
                                char22_2[49] <= 32'h00003F00;
                                char22_2[50] <= 32'h00003F00;
                                char22_2[51] <= 32'h00007F80;
                                char22_2[52] <= 32'h000FFFFC;
                                char22_2[53] <= 32'h000FFFFC;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//4
                            4'd5: begin
                                char22_2[  0] <= 32'h00000000;
                                char22_2[  1] <= 32'h00000000;
                                char22_2[  2] <= 32'h00000000;
                                char22_2[  3] <= 32'h00000000;
                                char22_2[  4] <= 32'h00000000;
                                char22_2[  5] <= 32'h00000000;
                                char22_2[  6] <= 32'h00000000;
                                char22_2[  7] <= 32'h00000000;
                                char22_2[  8] <= 32'h00000000;
                                char22_2[  9] <= 32'h00000000;
                                char22_2[10] <= 32'h00000000;
                                char22_2[11] <= 32'h03FFFFF0;
                                char22_2[12] <= 32'h03FFFFF0;
                                char22_2[13] <= 32'h03FFFFF0;
                                char22_2[14] <= 32'h03FFFFE0;
                                char22_2[15] <= 32'h03800000;
                                char22_2[16] <= 32'h03800000;
                                char22_2[17] <= 32'h03800000;
                                char22_2[18] <= 32'h03800000;
                                char22_2[19] <= 32'h03800000;
                                char22_2[20] <= 32'h07800000;
                                char22_2[21] <= 32'h07800000;
                                char22_2[22] <= 32'h07800000;
                                char22_2[23] <= 32'h07800000;
                                char22_2[24] <= 32'h07800000;
                                char22_2[25] <= 32'h07800000;
                                char22_2[26] <= 32'h078FF800;
                                char22_2[27] <= 32'h073FFE00;
                                char22_2[28] <= 32'h077FFF80;
                                char22_2[29] <= 32'h07FC3F80;
                                char22_2[30] <= 32'h07E00FC0;
                                char22_2[31] <= 32'h07C007E0;
                                char22_2[32] <= 32'h078007E0;
                                char22_2[33] <= 32'h078003F0;
                                char22_2[34] <= 32'h000003F0;
                                char22_2[35] <= 32'h000001F0;
                                char22_2[36] <= 32'h000001F8;
                                char22_2[37] <= 32'h000001F8;
                                char22_2[38] <= 32'h000001F8;
                                char22_2[39] <= 32'h000001F8;
                                char22_2[40] <= 32'h000001F8;
                                char22_2[41] <= 32'h078001F8;
                                char22_2[42] <= 32'h0FC001F8;
                                char22_2[43] <= 32'h1FC001F0;
                                char22_2[44] <= 32'h1FC001F0;
                                char22_2[45] <= 32'h1FC003F0;
                                char22_2[46] <= 32'h1F8003F0;
                                char22_2[47] <= 32'h1F8003E0;
                                char22_2[48] <= 32'h0F8007E0;
                                char22_2[49] <= 32'h078007C0;
                                char22_2[50] <= 32'h07C01F80;
                                char22_2[51] <= 32'h03F83F00;
                                char22_2[52] <= 32'h00FFFE00;
                                char22_2[53] <= 32'h003FF800;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//5
                            4'd6: begin
                                char22_2[0] <= 32'h00000000;
                                char22_2[1] <= 32'h00000000;
                                char22_2[2] <= 32'h00000000;
                                char22_2[3] <= 32'h00000000;
                                char22_2[4] <= 32'h00000000;
                                char22_2[5] <= 32'h00000000;
                                char22_2[6] <= 32'h00000000;
                                char22_2[7] <= 32'h00000000;
                                char22_2[8] <= 32'h00000000;
                                char22_2[9] <= 32'h00000000;
                                char22_2[10] <= 32'h0007FE00;
                                char22_2[11] <= 32'h001FFF80;
                                char22_2[12] <= 32'h003F0FC0;
                                char22_2[13] <= 32'h007C07C0;
                                char22_2[14] <= 32'h00F807E0;
                                char22_2[15] <= 32'h01F007E0;
                                char22_2[16] <= 32'h03E007E0;
                                char22_2[17] <= 32'h03C007E0;
                                char22_2[18] <= 32'h07C003C0;
                                char22_2[19] <= 32'h07C00000;
                                char22_2[20] <= 32'h0FC00000;
                                char22_2[21] <= 32'h0F800000;
                                char22_2[22] <= 32'h0F800000;
                                char22_2[23] <= 32'h1F800000;
                                char22_2[24] <= 32'h1F800000;
                                char22_2[25] <= 32'h1F800000;
                                char22_2[26] <= 32'h1F87FE00;
                                char22_2[27] <= 32'h1F9FFF80;
                                char22_2[28] <= 32'h1FBFFFC0;
                                char22_2[29] <= 32'h3FFE1FC0;
                                char22_2[30] <= 32'h3FF807E0;
                                char22_2[31] <= 32'h3FE003F0;
                                char22_2[32] <= 32'h3FE003F0;
                                char22_2[33] <= 32'h3FC001F8;
                                char22_2[34] <= 32'h3F8001F8;
                                char22_2[35] <= 32'h3F8001F8;
                                char22_2[36] <= 32'h3F8000F8;
                                char22_2[37] <= 32'h3F8000F8;
                                char22_2[38] <= 32'h3F8000F8;
                                char22_2[39] <= 32'h1F8000F8;
                                char22_2[40] <= 32'h1F8000F8;
                                char22_2[41] <= 32'h1F8000F8;
                                char22_2[42] <= 32'h1F8000F8;
                                char22_2[43] <= 32'h1F8000F8;
                                char22_2[44] <= 32'h0FC001F8;
                                char22_2[45] <= 32'h0FC001F8;
                                char22_2[46] <= 32'h0FC001F0;
                                char22_2[47] <= 32'h07E001F0;
                                char22_2[48] <= 32'h03E003E0;
                                char22_2[49] <= 32'h03F003E0;
                                char22_2[50] <= 32'h01F807C0;
                                char22_2[51] <= 32'h00FE1F80;
                                char22_2[52] <= 32'h007FFE00;
                                char22_2[53] <= 32'h001FF800;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//6
                            4'd7: begin
                                char22_2[0] <= 32'h00000000;
                                char22_2[1] <= 32'h00000000;
                                char22_2[2] <= 32'h00000000;
                                char22_2[3] <= 32'h00000000;
                                char22_2[4] <= 32'h00000000;
                                char22_2[5] <= 32'h00000000;
                                char22_2[6] <= 32'h00000000;
                                char22_2[7] <= 32'h00000000;
                                char22_2[8] <= 32'h00000000;
                                char22_2[9] <= 32'h00000000;
                                char22_2[10] <= 32'h00000000;
                                char22_2[11] <= 32'h07FFFFF8;
                                char22_2[12] <= 32'h07FFFFF8;
                                char22_2[13] <= 32'h07FFFFF8;
                                char22_2[14] <= 32'h0FFFFFF0;
                                char22_2[15] <= 32'h0FC000E0;
                                char22_2[16] <= 32'h0F8001E0;
                                char22_2[17] <= 32'h0F0001C0;
                                char22_2[18] <= 32'h0E0003C0;
                                char22_2[19] <= 32'h0E000780;
                                char22_2[20] <= 32'h1E000780;
                                char22_2[21] <= 32'h1C000F00;
                                char22_2[22] <= 32'h00000F00;
                                char22_2[23] <= 32'h00001E00;
                                char22_2[24] <= 32'h00001E00;
                                char22_2[25] <= 32'h00003C00;
                                char22_2[26] <= 32'h00003C00;
                                char22_2[27] <= 32'h00007800;
                                char22_2[28] <= 32'h00007800;
                                char22_2[29] <= 32'h0000F800;
                                char22_2[30] <= 32'h0000F000;
                                char22_2[31] <= 32'h0001F000;
                                char22_2[32] <= 32'h0001E000;
                                char22_2[33] <= 32'h0003E000;
                                char22_2[34] <= 32'h0003E000;
                                char22_2[35] <= 32'h0003E000;
                                char22_2[36] <= 32'h0007C000;
                                char22_2[37] <= 32'h0007C000;
                                char22_2[38] <= 32'h0007C000;
                                char22_2[39] <= 32'h000FC000;
                                char22_2[40] <= 32'h000FC000;
                                char22_2[41] <= 32'h000FC000;
                                char22_2[42] <= 32'h000FC000;
                                char22_2[43] <= 32'h001FC000;
                                char22_2[44] <= 32'h001FC000;
                                char22_2[45] <= 32'h001FC000;
                                char22_2[46] <= 32'h001FC000;
                                char22_2[47] <= 32'h001FC000;
                                char22_2[48] <= 32'h001FC000;
                                char22_2[49] <= 32'h001FC000;
                                char22_2[50] <= 32'h001FC000;
                                char22_2[51] <= 32'h001FC000;
                                char22_2[52] <= 32'h001FC000;
                                char22_2[53] <= 32'h000F8000;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//7
                            4'd8: begin
                                char22_2[0] <= 32'h00000000;
                                char22_2[1] <= 32'h00000000;
                                char22_2[2] <= 32'h00000000;
                                char22_2[3] <= 32'h00000000;
                                char22_2[4] <= 32'h00000000;
                                char22_2[5] <= 32'h00000000;
                                char22_2[6] <= 32'h00000000;
                                char22_2[7] <= 32'h00000000;
                                char22_2[8] <= 32'h00000000;
                                char22_2[9] <= 32'h00000000;
                                char22_2[10] <= 32'h003FF800;
                                char22_2[11] <= 32'h00FFFE00;
                                char22_2[12] <= 32'h01F81F80;
                                char22_2[13] <= 32'h03E00FC0;
                                char22_2[14] <= 32'h07C003E0;
                                char22_2[15] <= 32'h0F8003E0;
                                char22_2[16] <= 32'h0F8001F0;
                                char22_2[17] <= 32'h1F0001F0;
                                char22_2[18] <= 32'h1F0001F0;
                                char22_2[19] <= 32'h1F0001F0;
                                char22_2[20] <= 32'h1F0001F0;
                                char22_2[21] <= 32'h1F0001F0;
                                char22_2[22] <= 32'h1F8001F0;
                                char22_2[23] <= 32'h1FC001F0;
                                char22_2[24] <= 32'h0FC001F0;
                                char22_2[25] <= 32'h0FF003E0;
                                char22_2[26] <= 32'h07F803C0;
                                char22_2[27] <= 32'h03FE0F80;
                                char22_2[28] <= 32'h01FF9F00;
                                char22_2[29] <= 32'h00FFFE00;
                                char22_2[30] <= 32'h003FF800;
                                char22_2[31] <= 32'h007FFC00;
                                char22_2[32] <= 32'h01F7FF00;
                                char22_2[33] <= 32'h03E1FF80;
                                char22_2[34] <= 32'h07C07FC0;
                                char22_2[35] <= 32'h0F801FE0;
                                char22_2[36] <= 32'h0F800FE0;
                                char22_2[37] <= 32'h1F0007F0;
                                char22_2[38] <= 32'h1F0003F0;
                                char22_2[39] <= 32'h3E0001F8;
                                char22_2[40] <= 32'h3E0001F8;
                                char22_2[41] <= 32'h3E0001F8;
                                char22_2[42] <= 32'h3E0000F8;
                                char22_2[43] <= 32'h3E0000F8;
                                char22_2[44] <= 32'h3E0000F8;
                                char22_2[45] <= 32'h3E0000F8;
                                char22_2[46] <= 32'h1F0001F0;
                                char22_2[47] <= 32'h1F0001F0;
                                char22_2[48] <= 32'h0F8003E0;
                                char22_2[49] <= 32'h0FC003E0;
                                char22_2[50] <= 32'h07E007C0;
                                char22_2[51] <= 32'h01F83F80;
                                char22_2[52] <= 32'h00FFFE00;
                                char22_2[53] <= 32'h003FF800;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//8
                            4'd9: begin
                                char22_2[0] <= 32'h00000000;
                                char22_2[1] <= 32'h00000000;
                                char22_2[2] <= 32'h00000000;
                                char22_2[3] <= 32'h00000000;
                                char22_2[4] <= 32'h00000000;
                                char22_2[5] <= 32'h00000000;
                                char22_2[6] <= 32'h00000000;
                                char22_2[7] <= 32'h00000000;
                                char22_2[8] <= 32'h00000000;
                                char22_2[9] <= 32'h00000000;
                                char22_2[10] <= 32'h003FF000;
                                char22_2[11] <= 32'h00FFFC00;
                                char22_2[12] <= 32'h01F83F00;
                                char22_2[13] <= 32'h03E01F80;
                                char22_2[14] <= 32'h07C00F80;
                                char22_2[15] <= 32'h0FC007C0;
                                char22_2[16] <= 32'h0F8003E0;
                                char22_2[17] <= 32'h1F8003E0;
                                char22_2[18] <= 32'h1F0003F0;
                                char22_2[19] <= 32'h1F0003F0;
                                char22_2[20] <= 32'h3F0001F0;
                                char22_2[21] <= 32'h3F0001F0;
                                char22_2[22] <= 32'h3F0001F8;
                                char22_2[23] <= 32'h3F0001F8;
                                char22_2[24] <= 32'h3F0001F8;
                                char22_2[25] <= 32'h3F0001F8;
                                char22_2[26] <= 32'h3F0001F8;
                                char22_2[27] <= 32'h3F0001F8;
                                char22_2[28] <= 32'h3F0003F8;
                                char22_2[29] <= 32'h1F8003F8;
                                char22_2[30] <= 32'h1F8007F8;
                                char22_2[31] <= 32'h1F800FF8;
                                char22_2[32] <= 32'h0FC01FF8;
                                char22_2[33] <= 32'h0FE03FF8;
                                char22_2[34] <= 32'h07F8FDF8;
                                char22_2[35] <= 32'h03FFF9F8;
                                char22_2[36] <= 32'h01FFF1F8;
                                char22_2[37] <= 32'h003F83F8;
                                char22_2[38] <= 32'h000003F0;
                                char22_2[39] <= 32'h000003F0;
                                char22_2[40] <= 32'h000003F0;
                                char22_2[41] <= 32'h000003F0;
                                char22_2[42] <= 32'h000007E0;
                                char22_2[43] <= 32'h000007E0;
                                char22_2[44] <= 32'h000007C0;
                                char22_2[45] <= 32'h03C007C0;
                                char22_2[46] <= 32'h07C00F80;
                                char22_2[47] <= 32'h0FE00F80;
                                char22_2[48] <= 32'h0FE01F00;
                                char22_2[49] <= 32'h0FE03E00;
                                char22_2[50] <= 32'h07E07E00;
                                char22_2[51] <= 32'h07F1F800;
                                char22_2[52] <= 32'h03FFF000;
                                char22_2[53] <= 32'h00FFC000;
                                char22_2[54] <= 32'h00000000;
                                char22_2[55] <= 32'h00000000;
                                char22_2[56] <= 32'h00000000;
                                char22_2[57] <= 32'h00000000;
                                char22_2[58] <= 32'h00000000;
                                char22_2[59] <= 32'h00000000;
                                char22_2[60] <= 32'h00000000;
                                char22_2[61] <= 32'h00000000;
                                char22_2[62] <= 32'h00000000;
                                char22_2[63] <= 32'h00000000;
                            end//9
                            default: begin
                                char22_2[0] <= char22_2[0];
                                char22_2[1] <= char22_2[1];
                                char22_2[2] <= char22_2[2];
                                char22_2[3] <= char22_2[3];
                                char22_2[4] <= char22_2[4];
                                char22_2[5] <= char22_2[5];
                                char22_2[6] <= char22_2[6];
                                char22_2[7] <= char22_2[7];
                                char22_2[8] <= char22_2[8];
                                char22_2[9] <= char22_2[9];
                                char22_2[10] <= char22_2[10];
                                char22_2[11] <= char22_2[11];
                                char22_2[12] <= char22_2[12];
                                char22_2[13] <= char22_2[13];
                                char22_2[14] <= char22_2[14];
                                char22_2[15] <= char22_2[15];
                                char22_2[16] <= char22_2[16];
                                char22_2[17] <= char22_2[17];
                                char22_2[18] <= char22_2[18];
                                char22_2[19] <= char22_2[19];
                                char22_2[20] <= char22_2[20];
                                char22_2[21] <= char22_2[21];
                                char22_2[22] <= char22_2[22];
                                char22_2[23] <= char22_2[23];
                                char22_2[24] <= char22_2[24];
                                char22_2[25] <= char22_2[25];
                                char22_2[26] <= char22_2[26];
                                char22_2[27] <= char22_2[27];
                                char22_2[28] <= char22_2[28];
                                char22_2[29] <= char22_2[29];
                                char22_2[30] <= char22_2[30];
                                char22_2[31] <= char22_2[31];
                                char22_2[32] <= char22_2[32];
                                char22_2[33] <= char22_2[33];
                                char22_2[34] <= char22_2[34];
                                char22_2[35] <= char22_2[35];
                                char22_2[36] <= char22_2[36];
                                char22_2[37] <= char22_2[37];
                                char22_2[38] <= char22_2[38];
                                char22_2[39] <= char22_2[39];
                                char22_2[40] <= char22_2[40];
                                char22_2[41] <= char22_2[41];
                                char22_2[42] <= char22_2[42];
                                char22_2[43] <= char22_2[43];
                                char22_2[44] <= char22_2[44];
                                char22_2[45] <= char22_2[45];
                                char22_2[46] <= char22_2[46];
                                char22_2[47] <= char22_2[47];
                                char22_2[48] <= char22_2[48];
                                char22_2[49] <= char22_2[49];
                                char22_2[50] <= char22_2[50];
                                char22_2[51] <= char22_2[51];
                                char22_2[52] <= char22_2[52];
                                char22_2[53] <= char22_2[53];
                                char22_2[54] <= char22_2[54];
                                char22_2[55] <= char22_2[55];
                                char22_2[56] <= char22_2[56];
                                char22_2[57] <= char22_2[57];
                                char22_2[58] <= char22_2[58];
                                char22_2[59] <= char22_2[59];
                                char22_2[60] <= char22_2[60];
                                char22_2[61] <= char22_2[61];
                                char22_2[62] <= char22_2[62];
                                char22_2[63] <= char22_2[63];
                            end
                        endcase
            
                 case((a0 - h1*(a0/h1))/t1)
                                4'd0: begin
                                    char22_3[  0] <= 32'h00000000;
                                    char22_3[  1] <= 32'h00000000;
                                    char22_3[  2] <= 32'h00000000;
                                    char22_3[  3] <= 32'h00000000;
                                    char22_3[  4] <= 32'h00000000;
                                    char22_3[  5] <= 32'h00000000;
                                    char22_3[  6] <= 32'h00000000;
                                    char22_3[  7] <= 32'h00000000;
                                    char22_3[  8] <= 32'h00000000;
                                    char22_3[  9] <= 32'h00000000;
                                    char22_3[10] <= 32'h000FF000;
                                    char22_3[11] <= 32'h003FFC00;
                                    char22_3[12] <= 32'h007E7E00;
                                    char22_3[13] <= 32'h00F81F00;
                                    char22_3[14] <= 32'h01F00F80;
                                    char22_3[15] <= 32'h03F00FC0;
                                    char22_3[16] <= 32'h03E007C0;
                                    char22_3[17] <= 32'h07E007E0;
                                    char22_3[18] <= 32'h07C003E0;
                                    char22_3[19] <= 32'h0FC003F0;
                                    char22_3[20] <= 32'h0FC003F0;
                                    char22_3[21] <= 32'h0FC003F0;
                                    char22_3[22] <= 32'h1F8001F8;
                                    char22_3[23] <= 32'h1F8001F8;
                                    char22_3[24] <= 32'h1F8001F8;
                                    char22_3[25] <= 32'h1F8001F8;
                                    char22_3[26] <= 32'h1F8001F8;
                                    char22_3[27] <= 32'h3F8001F8;
                                    char22_3[28] <= 32'h3F8001F8;
                                    char22_3[29] <= 32'h3F8001F8;
                                    char22_3[30] <= 32'h3F8001F8;
                                    char22_3[31] <= 32'h3F8001F8;
                                    char22_3[32] <= 32'h3F8001F8;
                                    char22_3[33] <= 32'h3F8001F8;
                                    char22_3[34] <= 32'h3F8001F8;
                                    char22_3[35] <= 32'h3F8001F8;
                                    char22_3[36] <= 32'h3F8001F8;
                                    char22_3[37] <= 32'h1F8001F8;
                                    char22_3[38] <= 32'h1F8001F8;
                                    char22_3[39] <= 32'h1F8001F8;
                                    char22_3[40] <= 32'h1F8001F8;
                                    char22_3[41] <= 32'h1F8001F0;
                                    char22_3[42] <= 32'h0F8003F0;
                                    char22_3[43] <= 32'h0FC003F0;
                                    char22_3[44] <= 32'h0FC003F0;
                                    char22_3[45] <= 32'h07C003E0;
                                    char22_3[46] <= 32'h07E007E0;
                                    char22_3[47] <= 32'h03E007C0;
                                    char22_3[48] <= 32'h03F00FC0;
                                    char22_3[49] <= 32'h01F00F80;
                                    char22_3[50] <= 32'h00F81F00;
                                    char22_3[51] <= 32'h007E7E00;
                                    char22_3[52] <= 32'h003FFC00;
                                    char22_3[53] <= 32'h000FF000;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//0
                                4'd1: begin
                                    char22_3[  0] <= 32'h00000000;
                                    char22_3[  1] <= 32'h00000000;
                                    char22_3[  2] <= 32'h00000000;
                                    char22_3[  3] <= 32'h00000000;
                                    char22_3[  4] <= 32'h00000000;
                                    char22_3[  5] <= 32'h00000000;
                                    char22_3[  6] <= 32'h00000000;
                                    char22_3[  7] <= 32'h00000000;
                                    char22_3[  8] <= 32'h00000000;
                                    char22_3[  9] <= 32'h00000000;
                                    char22_3[10] <= 32'h0000E000;
                                    char22_3[11] <= 32'h0001E000;
                                    char22_3[12] <= 32'h0003E000;
                                    char22_3[13] <= 32'h001FE000;
                                    char22_3[14] <= 32'h03FFE000;
                                    char22_3[15] <= 32'h03FFE000;
                                    char22_3[16] <= 32'h0007E000;
                                    char22_3[17] <= 32'h0007E000;
                                    char22_3[18] <= 32'h0007E000;
                                    char22_3[19] <= 32'h0007E000;
                                    char22_3[20] <= 32'h0007E000;
                                    char22_3[21] <= 32'h0007E000;
                                    char22_3[22] <= 32'h0007E000;
                                    char22_3[23] <= 32'h0007E000;
                                    char22_3[24] <= 32'h0007E000;
                                    char22_3[25] <= 32'h0007E000;
                                    char22_3[26] <= 32'h0007E000;
                                    char22_3[27] <= 32'h0007E000;
                                    char22_3[28] <= 32'h0007E000;
                                    char22_3[29] <= 32'h0007E000;
                                    char22_3[30] <= 32'h0007E000;
                                    char22_3[31] <= 32'h0007E000;
                                    char22_3[32] <= 32'h0007E000;
                                    char22_3[33] <= 32'h0007E000;
                                    char22_3[34] <= 32'h0007E000;
                                    char22_3[35] <= 32'h0007E000;
                                    char22_3[36] <= 32'h0007E000;
                                    char22_3[37] <= 32'h0007E000;
                                    char22_3[38] <= 32'h0007E000;
                                    char22_3[39] <= 32'h0007E000;
                                    char22_3[40] <= 32'h0007E000;
                                    char22_3[41] <= 32'h0007E000;
                                    char22_3[42] <= 32'h0007E000;
                                    char22_3[43] <= 32'h0007E000;
                                    char22_3[44] <= 32'h0007E000;
                                    char22_3[45] <= 32'h0007E000;
                                    char22_3[46] <= 32'h0007E000;
                                    char22_3[47] <= 32'h0007E000;
                                    char22_3[48] <= 32'h0007E000;
                                    char22_3[49] <= 32'h0007E000;
                                    char22_3[50] <= 32'h0007E000;
                                    char22_3[51] <= 32'h000FF800;
                                    char22_3[52] <= 32'h03FFFFC0;
                                    char22_3[53] <= 32'h03FFFFC0;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//1
                                4'd2: begin
                                    char22_3[  0] <= 32'h00000000;
                                    char22_3[  1] <= 32'h00000000;
                                    char22_3[  2] <= 32'h00000000;
                                    char22_3[  3] <= 32'h00000000;
                                    char22_3[  4] <= 32'h00000000;
                                    char22_3[  5] <= 32'h00000000;
                                    char22_3[  6] <= 32'h00000000;
                                    char22_3[  7] <= 32'h00000000;
                                    char22_3[  8] <= 32'h00000000;
                                    char22_3[  9] <= 32'h00000000;
                                    char22_3[10] <= 32'h001FFC00;
                                    char22_3[11] <= 32'h007FFF00;
                                    char22_3[12] <= 32'h01F83F80;
                                    char22_3[13] <= 32'h03E00FC0;
                                    char22_3[14] <= 32'h07C007E0;
                                    char22_3[15] <= 32'h078007E0;
                                    char22_3[16] <= 32'h0F8003F0;
                                    char22_3[17] <= 32'h0F8003F0;
                                    char22_3[18] <= 32'h1F8003F0;
                                    char22_3[19] <= 32'h1F8003F0;
                                    char22_3[20] <= 32'h1FC003F0;
                                    char22_3[21] <= 32'h1FC003F0;
                                    char22_3[22] <= 32'h1FC003F0;
                                    char22_3[23] <= 32'h0FC003F0;
                                    char22_3[24] <= 32'h07C003F0;
                                    char22_3[25] <= 32'h000003E0;
                                    char22_3[26] <= 32'h000007E0;
                                    char22_3[27] <= 32'h000007E0;
                                    char22_3[28] <= 32'h00000FC0;
                                    char22_3[29] <= 32'h00000F80;
                                    char22_3[30] <= 32'h00001F80;
                                    char22_3[31] <= 32'h00003F00;
                                    char22_3[32] <= 32'h00003E00;
                                    char22_3[33] <= 32'h00007C00;
                                    char22_3[34] <= 32'h0000F800;
                                    char22_3[35] <= 32'h0001F000;
                                    char22_3[36] <= 32'h0003E000;
                                    char22_3[37] <= 32'h0007C000;
                                    char22_3[38] <= 32'h000F8000;
                                    char22_3[39] <= 32'h001F0000;
                                    char22_3[40] <= 32'h003E0000;
                                    char22_3[41] <= 32'h007C0000;
                                    char22_3[42] <= 32'h00F80000;
                                    char22_3[43] <= 32'h01F00038;
                                    char22_3[44] <= 32'h01E00038;
                                    char22_3[45] <= 32'h03C00070;
                                    char22_3[46] <= 32'h07800070;
                                    char22_3[47] <= 32'h0F8000F0;
                                    char22_3[48] <= 32'h0F0000F0;
                                    char22_3[49] <= 32'h1E0003F0;
                                    char22_3[50] <= 32'h3FFFFFF0;
                                    char22_3[51] <= 32'h3FFFFFF0;
                                    char22_3[52] <= 32'h3FFFFFE0;
                                    char22_3[53] <= 32'h3FFFFFE0;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//2
                                4'd3: begin
                                    char22_3[  0] <= 32'h00000000;
                                    char22_3[  1] <= 32'h00000000;
                                    char22_3[  2] <= 32'h00000000;
                                    char22_3[  3] <= 32'h00000000;
                                    char22_3[  4] <= 32'h00000000;
                                    char22_3[  5] <= 32'h00000000;
                                    char22_3[  6] <= 32'h00000000;
                                    char22_3[  7] <= 32'h00000000;
                                    char22_3[  8] <= 32'h00000000;
                                    char22_3[  9] <= 32'h00000000;
                                    char22_3[10] <= 32'h003FF000;
                                    char22_3[11] <= 32'h00FFFC00;
                                    char22_3[12] <= 32'h01F07E00;
                                    char22_3[13] <= 32'h03C03F00;
                                    char22_3[14] <= 32'h07801F80;
                                    char22_3[15] <= 32'h0F800FC0;
                                    char22_3[16] <= 32'h0F800FC0;
                                    char22_3[17] <= 32'h0F8007E0;
                                    char22_3[18] <= 32'h0FC007E0;
                                    char22_3[19] <= 32'h0FC007E0;
                                    char22_3[20] <= 32'h0FC007E0;
                                    char22_3[21] <= 32'h07C007E0;
                                    char22_3[22] <= 32'h000007E0;
                                    char22_3[23] <= 32'h000007E0;
                                    char22_3[24] <= 32'h000007C0;
                                    char22_3[25] <= 32'h00000FC0;
                                    char22_3[26] <= 32'h00000F80;
                                    char22_3[27] <= 32'h00001F00;
                                    char22_3[28] <= 32'h00007E00;
                                    char22_3[29] <= 32'h0003FC00;
                                    char22_3[30] <= 32'h001FF000;
                                    char22_3[31] <= 32'h001FFC00;
                                    char22_3[32] <= 32'h0000FF00;
                                    char22_3[33] <= 32'h00001F80;
                                    char22_3[34] <= 32'h00000FC0;
                                    char22_3[35] <= 32'h000007E0;
                                    char22_3[36] <= 32'h000003E0;
                                    char22_3[37] <= 32'h000003F0;
                                    char22_3[38] <= 32'h000003F0;
                                    char22_3[39] <= 32'h000001F0;
                                    char22_3[40] <= 32'h000001F8;
                                    char22_3[41] <= 32'h000001F8;
                                    char22_3[42] <= 32'h078001F8;
                                    char22_3[43] <= 32'h0FC001F8;
                                    char22_3[44] <= 32'h1FC001F8;
                                    char22_3[45] <= 32'h1FC003F0;
                                    char22_3[46] <= 32'h1FC003F0;
                                    char22_3[47] <= 32'h1FC003E0;
                                    char22_3[48] <= 32'h0F8007E0;
                                    char22_3[49] <= 32'h0F8007C0;
                                    char22_3[50] <= 32'h07C01F80;
                                    char22_3[51] <= 32'h03F07F00;
                                    char22_3[52] <= 32'h01FFFE00;
                                    char22_3[53] <= 32'h003FF000;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//3
                                4'd4: begin
                                    char22_3[  0] <= 32'h00000000;
                                    char22_3[  1] <= 32'h00000000;
                                    char22_3[  2] <= 32'h00000000;
                                    char22_3[  3] <= 32'h00000000;
                                    char22_3[  4] <= 32'h00000000;
                                    char22_3[  5] <= 32'h00000000;
                                    char22_3[  6] <= 32'h00000000;
                                    char22_3[  7] <= 32'h00000000;
                                    char22_3[  8] <= 32'h00000000;
                                    char22_3[  9] <= 32'h00000000;
                                    char22_3[10] <= 32'h00001F00;
                                    char22_3[11] <= 32'h00001F00;
                                    char22_3[12] <= 32'h00003F00;
                                    char22_3[13] <= 32'h00003F00;
                                    char22_3[14] <= 32'h00007F00;
                                    char22_3[15] <= 32'h0000FF00;
                                    char22_3[16] <= 32'h0000FF00;
                                    char22_3[17] <= 32'h0001FF00;
                                    char22_3[18] <= 32'h0003FF00;
                                    char22_3[19] <= 32'h0003BF00;
                                    char22_3[20] <= 32'h0007BF00;
                                    char22_3[21] <= 32'h00073F00;
                                    char22_3[22] <= 32'h000F3F00;
                                    char22_3[23] <= 32'h001E3F00;
                                    char22_3[24] <= 32'h001C3F00;
                                    char22_3[25] <= 32'h003C3F00;
                                    char22_3[26] <= 32'h00783F00;
                                    char22_3[27] <= 32'h00783F00;
                                    char22_3[28] <= 32'h00F03F00;
                                    char22_3[29] <= 32'h00E03F00;
                                    char22_3[30] <= 32'h01E03F00;
                                    char22_3[31] <= 32'h03C03F00;
                                    char22_3[32] <= 32'h03803F00;
                                    char22_3[33] <= 32'h07803F00;
                                    char22_3[34] <= 32'h0F003F00;
                                    char22_3[35] <= 32'h0F003F00;
                                    char22_3[36] <= 32'h1E003F00;
                                    char22_3[37] <= 32'h1C003F00;
                                    char22_3[38] <= 32'h3C003F00;
                                    char22_3[39] <= 32'h7FFFFFFE;
                                    char22_3[40] <= 32'h7FFFFFFE;
                                    char22_3[41] <= 32'h00003F00;
                                    char22_3[42] <= 32'h00003F00;
                                    char22_3[43] <= 32'h00003F00;
                                    char22_3[44] <= 32'h00003F00;
                                    char22_3[45] <= 32'h00003F00;
                                    char22_3[46] <= 32'h00003F00;
                                    char22_3[47] <= 32'h00003F00;
                                    char22_3[48] <= 32'h00003F00;
                                    char22_3[49] <= 32'h00003F00;
                                    char22_3[50] <= 32'h00003F00;
                                    char22_3[51] <= 32'h00007F80;
                                    char22_3[52] <= 32'h000FFFFC;
                                    char22_3[53] <= 32'h000FFFFC;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//4
                                4'd5: begin
                                    char22_3[  0] <= 32'h00000000;
                                    char22_3[  1] <= 32'h00000000;
                                    char22_3[  2] <= 32'h00000000;
                                    char22_3[  3] <= 32'h00000000;
                                    char22_3[  4] <= 32'h00000000;
                                    char22_3[  5] <= 32'h00000000;
                                    char22_3[  6] <= 32'h00000000;
                                    char22_3[  7] <= 32'h00000000;
                                    char22_3[  8] <= 32'h00000000;
                                    char22_3[  9] <= 32'h00000000;
                                    char22_3[10] <= 32'h00000000;
                                    char22_3[11] <= 32'h03FFFFF0;
                                    char22_3[12] <= 32'h03FFFFF0;
                                    char22_3[13] <= 32'h03FFFFF0;
                                    char22_3[14] <= 32'h03FFFFE0;
                                    char22_3[15] <= 32'h03800000;
                                    char22_3[16] <= 32'h03800000;
                                    char22_3[17] <= 32'h03800000;
                                    char22_3[18] <= 32'h03800000;
                                    char22_3[19] <= 32'h03800000;
                                    char22_3[20] <= 32'h07800000;
                                    char22_3[21] <= 32'h07800000;
                                    char22_3[22] <= 32'h07800000;
                                    char22_3[23] <= 32'h07800000;
                                    char22_3[24] <= 32'h07800000;
                                    char22_3[25] <= 32'h07800000;
                                    char22_3[26] <= 32'h078FF800;
                                    char22_3[27] <= 32'h073FFE00;
                                    char22_3[28] <= 32'h077FFF80;
                                    char22_3[29] <= 32'h07FC3F80;
                                    char22_3[30] <= 32'h07E00FC0;
                                    char22_3[31] <= 32'h07C007E0;
                                    char22_3[32] <= 32'h078007E0;
                                    char22_3[33] <= 32'h078003F0;
                                    char22_3[34] <= 32'h000003F0;
                                    char22_3[35] <= 32'h000001F0;
                                    char22_3[36] <= 32'h000001F8;
                                    char22_3[37] <= 32'h000001F8;
                                    char22_3[38] <= 32'h000001F8;
                                    char22_3[39] <= 32'h000001F8;
                                    char22_3[40] <= 32'h000001F8;
                                    char22_3[41] <= 32'h078001F8;
                                    char22_3[42] <= 32'h0FC001F8;
                                    char22_3[43] <= 32'h1FC001F0;
                                    char22_3[44] <= 32'h1FC001F0;
                                    char22_3[45] <= 32'h1FC003F0;
                                    char22_3[46] <= 32'h1F8003F0;
                                    char22_3[47] <= 32'h1F8003E0;
                                    char22_3[48] <= 32'h0F8007E0;
                                    char22_3[49] <= 32'h078007C0;
                                    char22_3[50] <= 32'h07C01F80;
                                    char22_3[51] <= 32'h03F83F00;
                                    char22_3[52] <= 32'h00FFFE00;
                                    char22_3[53] <= 32'h003FF800;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//5
                                4'd6: begin
                                    char22_3[0] <= 32'h00000000;
                                    char22_3[1] <= 32'h00000000;
                                    char22_3[2] <= 32'h00000000;
                                    char22_3[3] <= 32'h00000000;
                                    char22_3[4] <= 32'h00000000;
                                    char22_3[5] <= 32'h00000000;
                                    char22_3[6] <= 32'h00000000;
                                    char22_3[7] <= 32'h00000000;
                                    char22_3[8] <= 32'h00000000;
                                    char22_3[9] <= 32'h00000000;
                                    char22_3[10] <= 32'h0007FE00;
                                    char22_3[11] <= 32'h001FFF80;
                                    char22_3[12] <= 32'h003F0FC0;
                                    char22_3[13] <= 32'h007C07C0;
                                    char22_3[14] <= 32'h00F807E0;
                                    char22_3[15] <= 32'h01F007E0;
                                    char22_3[16] <= 32'h03E007E0;
                                    char22_3[17] <= 32'h03C007E0;
                                    char22_3[18] <= 32'h07C003C0;
                                    char22_3[19] <= 32'h07C00000;
                                    char22_3[20] <= 32'h0FC00000;
                                    char22_3[21] <= 32'h0F800000;
                                    char22_3[22] <= 32'h0F800000;
                                    char22_3[23] <= 32'h1F800000;
                                    char22_3[24] <= 32'h1F800000;
                                    char22_3[25] <= 32'h1F800000;
                                    char22_3[26] <= 32'h1F87FE00;
                                    char22_3[27] <= 32'h1F9FFF80;
                                    char22_3[28] <= 32'h1FBFFFC0;
                                    char22_3[29] <= 32'h3FFE1FC0;
                                    char22_3[30] <= 32'h3FF807E0;
                                    char22_3[31] <= 32'h3FE003F0;
                                    char22_3[32] <= 32'h3FE003F0;
                                    char22_3[33] <= 32'h3FC001F8;
                                    char22_3[34] <= 32'h3F8001F8;
                                    char22_3[35] <= 32'h3F8001F8;
                                    char22_3[36] <= 32'h3F8000F8;
                                    char22_3[37] <= 32'h3F8000F8;
                                    char22_3[38] <= 32'h3F8000F8;
                                    char22_3[39] <= 32'h1F8000F8;
                                    char22_3[40] <= 32'h1F8000F8;
                                    char22_3[41] <= 32'h1F8000F8;
                                    char22_3[42] <= 32'h1F8000F8;
                                    char22_3[43] <= 32'h1F8000F8;
                                    char22_3[44] <= 32'h0FC001F8;
                                    char22_3[45] <= 32'h0FC001F8;
                                    char22_3[46] <= 32'h0FC001F0;
                                    char22_3[47] <= 32'h07E001F0;
                                    char22_3[48] <= 32'h03E003E0;
                                    char22_3[49] <= 32'h03F003E0;
                                    char22_3[50] <= 32'h01F807C0;
                                    char22_3[51] <= 32'h00FE1F80;
                                    char22_3[52] <= 32'h007FFE00;
                                    char22_3[53] <= 32'h001FF800;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//6
                                4'd7: begin
                                    char22_3[0] <= 32'h00000000;
                                    char22_3[1] <= 32'h00000000;
                                    char22_3[2] <= 32'h00000000;
                                    char22_3[3] <= 32'h00000000;
                                    char22_3[4] <= 32'h00000000;
                                    char22_3[5] <= 32'h00000000;
                                    char22_3[6] <= 32'h00000000;
                                    char22_3[7] <= 32'h00000000;
                                    char22_3[8] <= 32'h00000000;
                                    char22_3[9] <= 32'h00000000;
                                    char22_3[10] <= 32'h00000000;
                                    char22_3[11] <= 32'h07FFFFF8;
                                    char22_3[12] <= 32'h07FFFFF8;
                                    char22_3[13] <= 32'h07FFFFF8;
                                    char22_3[14] <= 32'h0FFFFFF0;
                                    char22_3[15] <= 32'h0FC000E0;
                                    char22_3[16] <= 32'h0F8001E0;
                                    char22_3[17] <= 32'h0F0001C0;
                                    char22_3[18] <= 32'h0E0003C0;
                                    char22_3[19] <= 32'h0E000780;
                                    char22_3[20] <= 32'h1E000780;
                                    char22_3[21] <= 32'h1C000F00;
                                    char22_3[22] <= 32'h00000F00;
                                    char22_3[23] <= 32'h00001E00;
                                    char22_3[24] <= 32'h00001E00;
                                    char22_3[25] <= 32'h00003C00;
                                    char22_3[26] <= 32'h00003C00;
                                    char22_3[27] <= 32'h00007800;
                                    char22_3[28] <= 32'h00007800;
                                    char22_3[29] <= 32'h0000F800;
                                    char22_3[30] <= 32'h0000F000;
                                    char22_3[31] <= 32'h0001F000;
                                    char22_3[32] <= 32'h0001E000;
                                    char22_3[33] <= 32'h0003E000;
                                    char22_3[34] <= 32'h0003E000;
                                    char22_3[35] <= 32'h0003E000;
                                    char22_3[36] <= 32'h0007C000;
                                    char22_3[37] <= 32'h0007C000;
                                    char22_3[38] <= 32'h0007C000;
                                    char22_3[39] <= 32'h000FC000;
                                    char22_3[40] <= 32'h000FC000;
                                    char22_3[41] <= 32'h000FC000;
                                    char22_3[42] <= 32'h000FC000;
                                    char22_3[43] <= 32'h001FC000;
                                    char22_3[44] <= 32'h001FC000;
                                    char22_3[45] <= 32'h001FC000;
                                    char22_3[46] <= 32'h001FC000;
                                    char22_3[47] <= 32'h001FC000;
                                    char22_3[48] <= 32'h001FC000;
                                    char22_3[49] <= 32'h001FC000;
                                    char22_3[50] <= 32'h001FC000;
                                    char22_3[51] <= 32'h001FC000;
                                    char22_3[52] <= 32'h001FC000;
                                    char22_3[53] <= 32'h000F8000;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//7
                                4'd8: begin
                                    char22_3[0] <= 32'h00000000;
                                    char22_3[1] <= 32'h00000000;
                                    char22_3[2] <= 32'h00000000;
                                    char22_3[3] <= 32'h00000000;
                                    char22_3[4] <= 32'h00000000;
                                    char22_3[5] <= 32'h00000000;
                                    char22_3[6] <= 32'h00000000;
                                    char22_3[7] <= 32'h00000000;
                                    char22_3[8] <= 32'h00000000;
                                    char22_3[9] <= 32'h00000000;
                                    char22_3[10] <= 32'h003FF800;
                                    char22_3[11] <= 32'h00FFFE00;
                                    char22_3[12] <= 32'h01F81F80;
                                    char22_3[13] <= 32'h03E00FC0;
                                    char22_3[14] <= 32'h07C003E0;
                                    char22_3[15] <= 32'h0F8003E0;
                                    char22_3[16] <= 32'h0F8001F0;
                                    char22_3[17] <= 32'h1F0001F0;
                                    char22_3[18] <= 32'h1F0001F0;
                                    char22_3[19] <= 32'h1F0001F0;
                                    char22_3[20] <= 32'h1F0001F0;
                                    char22_3[21] <= 32'h1F0001F0;
                                    char22_3[22] <= 32'h1F8001F0;
                                    char22_3[23] <= 32'h1FC001F0;
                                    char22_3[24] <= 32'h0FC001F0;
                                    char22_3[25] <= 32'h0FF003E0;
                                    char22_3[26] <= 32'h07F803C0;
                                    char22_3[27] <= 32'h03FE0F80;
                                    char22_3[28] <= 32'h01FF9F00;
                                    char22_3[29] <= 32'h00FFFE00;
                                    char22_3[30] <= 32'h003FF800;
                                    char22_3[31] <= 32'h007FFC00;
                                    char22_3[32] <= 32'h01F7FF00;
                                    char22_3[33] <= 32'h03E1FF80;
                                    char22_3[34] <= 32'h07C07FC0;
                                    char22_3[35] <= 32'h0F801FE0;
                                    char22_3[36] <= 32'h0F800FE0;
                                    char22_3[37] <= 32'h1F0007F0;
                                    char22_3[38] <= 32'h1F0003F0;
                                    char22_3[39] <= 32'h3E0001F8;
                                    char22_3[40] <= 32'h3E0001F8;
                                    char22_3[41] <= 32'h3E0001F8;
                                    char22_3[42] <= 32'h3E0000F8;
                                    char22_3[43] <= 32'h3E0000F8;
                                    char22_3[44] <= 32'h3E0000F8;
                                    char22_3[45] <= 32'h3E0000F8;
                                    char22_3[46] <= 32'h1F0001F0;
                                    char22_3[47] <= 32'h1F0001F0;
                                    char22_3[48] <= 32'h0F8003E0;
                                    char22_3[49] <= 32'h0FC003E0;
                                    char22_3[50] <= 32'h07E007C0;
                                    char22_3[51] <= 32'h01F83F80;
                                    char22_3[52] <= 32'h00FFFE00;
                                    char22_3[53] <= 32'h003FF800;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//8
                                4'd9: begin
                                    char22_3[0] <= 32'h00000000;
                                    char22_3[1] <= 32'h00000000;
                                    char22_3[2] <= 32'h00000000;
                                    char22_3[3] <= 32'h00000000;
                                    char22_3[4] <= 32'h00000000;
                                    char22_3[5] <= 32'h00000000;
                                    char22_3[6] <= 32'h00000000;
                                    char22_3[7] <= 32'h00000000;
                                    char22_3[8] <= 32'h00000000;
                                    char22_3[9] <= 32'h00000000;
                                    char22_3[10] <= 32'h003FF000;
                                    char22_3[11] <= 32'h00FFFC00;
                                    char22_3[12] <= 32'h01F83F00;
                                    char22_3[13] <= 32'h03E01F80;
                                    char22_3[14] <= 32'h07C00F80;
                                    char22_3[15] <= 32'h0FC007C0;
                                    char22_3[16] <= 32'h0F8003E0;
                                    char22_3[17] <= 32'h1F8003E0;
                                    char22_3[18] <= 32'h1F0003F0;
                                    char22_3[19] <= 32'h1F0003F0;
                                    char22_3[20] <= 32'h3F0001F0;
                                    char22_3[21] <= 32'h3F0001F0;
                                    char22_3[22] <= 32'h3F0001F8;
                                    char22_3[23] <= 32'h3F0001F8;
                                    char22_3[24] <= 32'h3F0001F8;
                                    char22_3[25] <= 32'h3F0001F8;
                                    char22_3[26] <= 32'h3F0001F8;
                                    char22_3[27] <= 32'h3F0001F8;
                                    char22_3[28] <= 32'h3F0003F8;
                                    char22_3[29] <= 32'h1F8003F8;
                                    char22_3[30] <= 32'h1F8007F8;
                                    char22_3[31] <= 32'h1F800FF8;
                                    char22_3[32] <= 32'h0FC01FF8;
                                    char22_3[33] <= 32'h0FE03FF8;
                                    char22_3[34] <= 32'h07F8FDF8;
                                    char22_3[35] <= 32'h03FFF9F8;
                                    char22_3[36] <= 32'h01FFF1F8;
                                    char22_3[37] <= 32'h003F83F8;
                                    char22_3[38] <= 32'h000003F0;
                                    char22_3[39] <= 32'h000003F0;
                                    char22_3[40] <= 32'h000003F0;
                                    char22_3[41] <= 32'h000003F0;
                                    char22_3[42] <= 32'h000007E0;
                                    char22_3[43] <= 32'h000007E0;
                                    char22_3[44] <= 32'h000007C0;
                                    char22_3[45] <= 32'h03C007C0;
                                    char22_3[46] <= 32'h07C00F80;
                                    char22_3[47] <= 32'h0FE00F80;
                                    char22_3[48] <= 32'h0FE01F00;
                                    char22_3[49] <= 32'h0FE03E00;
                                    char22_3[50] <= 32'h07E07E00;
                                    char22_3[51] <= 32'h07F1F800;
                                    char22_3[52] <= 32'h03FFF000;
                                    char22_3[53] <= 32'h00FFC000;
                                    char22_3[54] <= 32'h00000000;
                                    char22_3[55] <= 32'h00000000;
                                    char22_3[56] <= 32'h00000000;
                                    char22_3[57] <= 32'h00000000;
                                    char22_3[58] <= 32'h00000000;
                                    char22_3[59] <= 32'h00000000;
                                    char22_3[60] <= 32'h00000000;
                                    char22_3[61] <= 32'h00000000;
                                    char22_3[62] <= 32'h00000000;
                                    char22_3[63] <= 32'h00000000;
                                end//9
                                default: begin
                                    char22_3[0] <= char22_3[0];
                                    char22_3[1] <= char22_3[1];
                                    char22_3[2] <= char22_3[2];
                                    char22_3[3] <= char22_3[3];
                                    char22_3[4] <= char22_3[4];
                                    char22_3[5] <= char22_3[5];
                                    char22_3[6] <= char22_3[6];
                                    char22_3[7] <= char22_3[7];
                                    char22_3[8] <= char22_3[8];
                                    char22_3[9] <= char22_3[9];
                                    char22_3[10] <= char22_3[10];
                                    char22_3[11] <= char22_3[11];
                                    char22_3[12] <= char22_3[12];
                                    char22_3[13] <= char22_3[13];
                                    char22_3[14] <= char22_3[14];
                                    char22_3[15] <= char22_3[15];
                                    char22_3[16] <= char22_3[16];
                                    char22_3[17] <= char22_3[17];
                                    char22_3[18] <= char22_3[18];
                                    char22_3[19] <= char22_3[19];
                                    char22_3[20] <= char22_3[20];
                                    char22_3[21] <= char22_3[21];
                                    char22_3[22] <= char22_3[22];
                                    char22_3[23] <= char22_3[23];
                                    char22_3[24] <= char22_3[24];
                                    char22_3[25] <= char22_3[25];
                                    char22_3[26] <= char22_3[26];
                                    char22_3[27] <= char22_3[27];
                                    char22_3[28] <= char22_3[28];
                                    char22_3[29] <= char22_3[29];
                                    char22_3[30] <= char22_3[30];
                                    char22_3[31] <= char22_3[31];
                                    char22_3[32] <= char22_3[32];
                                    char22_3[33] <= char22_3[33];
                                    char22_3[34] <= char22_3[34];
                                    char22_3[35] <= char22_3[35];
                                    char22_3[36] <= char22_3[36];
                                    char22_3[37] <= char22_3[37];
                                    char22_3[38] <= char22_3[38];
                                    char22_3[39] <= char22_3[39];
                                    char22_3[40] <= char22_3[40];
                                    char22_3[41] <= char22_3[41];
                                    char22_3[42] <= char22_3[42];
                                    char22_3[43] <= char22_3[43];
                                    char22_3[44] <= char22_3[44];
                                    char22_3[45] <= char22_3[45];
                                    char22_3[46] <= char22_3[46];
                                    char22_3[47] <= char22_3[47];
                                    char22_3[48] <= char22_3[48];
                                    char22_3[49] <= char22_3[49];
                                    char22_3[50] <= char22_3[50];
                                    char22_3[51] <= char22_3[51];
                                    char22_3[52] <= char22_3[52];
                                    char22_3[53] <= char22_3[53];
                                    char22_3[54] <= char22_3[54];
                                    char22_3[55] <= char22_3[55];
                                    char22_3[56] <= char22_3[56];
                                    char22_3[57] <= char22_3[57];
                                    char22_3[58] <= char22_3[58];
                                    char22_3[59] <= char22_3[59];
                                    char22_3[60] <= char22_3[60];
                                    char22_3[61] <= char22_3[61];
                                    char22_3[62] <= char22_3[62];
                                    char22_3[63] <= char22_3[63];
                                end
                            endcase
           
                case((a0 - t1*(a0/t1))/o1)
                           4'd0: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h000FF000000000000000000000000000;
                                 char22_4[11] <= 128'h003FFC00000000000000000000000000;
                                 char22_4[12] <= 128'h007E7E00800000000000000000000000;
                                 char22_4[13] <= 128'h00F81F00000000000000000000000000;
                                 char22_4[14] <= 128'h01F00F80000000000000000000000000;
                                 char22_4[15] <= 128'h03F00FC0000000000000000000000000;
                                 char22_4[16] <= 128'h03E007C0000000000000000000000000;
                                 char22_4[17] <= 128'h07E007E0000000000000000000000000;
                                 char22_4[18] <= 128'h07C003E0000000000000000000000000;
                                 char22_4[19] <= 128'h0FC003F0000000000000000000000000;
                                 char22_4[20] <= 128'h0FC003F0000000000000000000000000;
                                 char22_4[21] <= 128'h0FC003F0000000000000000000000000;
                                 char22_4[22] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[23] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[24] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[25] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[26] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[27] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[28] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[29] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[30] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[31] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[32] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[33] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[34] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[35] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[36] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[37] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[38] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[39] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[40] <= 128'h1F8001F8000000000000000000000000;
                                 char22_4[41] <= 128'h1F8001F0000000000000000000000000;
                                 char22_4[42] <= 128'h0F8003F0000000000000000000000000;
                                 char22_4[43] <= 128'h0FC003F0000000000000000000000000;
                                 char22_4[44] <= 128'h0FC003F0000000000000000000000000;
                                 char22_4[45] <= 128'h07C003E0000000000000000000000000;
                                 char22_4[46] <= 128'h07E007E0000000000000000000000000;
                                 char22_4[47] <= 128'h03E007C0000000000000000000000000;
                                 char22_4[48] <= 128'h03F00FC0000000000000000000000000;
                                 char22_4[49] <= 128'h01F00F80000000000000000000000000;
                                 char22_4[50] <= 128'h00F81F00000000000000000000000000;
                                 char22_4[51] <= 128'h007E7E00000000000000000000000000;
                                 char22_4[52] <= 128'h003FFC00000000000000000000000000;
                                 char22_4[53] <= 128'h000FF000000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//0
                           4'd1: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h0000E000000000000000000000000000;
                                 char22_4[11] <= 128'h0001E000000000000000000000000000;
                                 char22_4[12] <= 128'h0003E000000000000000000000000000;
                                 char22_4[13] <= 128'h001FE000000000000000000000000000;
                                 char22_4[14] <= 128'h03FFE000000000000000000000000000;
                                 char22_4[15] <= 128'h03FFE000000000000000000000000000;
                                 char22_4[16] <= 128'h0007E000000000000000000000000000;
                                 char22_4[17] <= 128'h0007E000000000000000000000000000;
                                 char22_4[18] <= 128'h0007E000000000000000000000000000;
                                 char22_4[19] <= 128'h0007E000000000000000000000000000;
                                 char22_4[20] <= 128'h0007E000000000000000000000000000;
                                 char22_4[21] <= 128'h0007E000000000000000000000000000;
                                 char22_4[22] <= 128'h0007E000000000000000000000000000;
                                 char22_4[23] <= 128'h0007E000000000000000000000000000;
                                 char22_4[24] <= 128'h0007E000000000000000000000000000;
                                 char22_4[25] <= 128'h0007E000000000000000000000000000;
                                 char22_4[26] <= 128'h0007E000000000000000000000000000;
                                 char22_4[27] <= 128'h0007E000000000000000000000000000;
                                 char22_4[28] <= 128'h0007E000000000000000000000000000;
                                 char22_4[29] <= 128'h0007E000000000000000000000000000;
                                 char22_4[30] <= 128'h0007E000000000000000000000000000;
                                 char22_4[31] <= 128'h0007E000000000000000000000000000;
                                 char22_4[32] <= 128'h0007E000000000000000000000000000;
                                 char22_4[33] <= 128'h0007E000000000000000000000000000;
                                 char22_4[34] <= 128'h0007E000000000000000000000000000;
                                 char22_4[35] <= 128'h0007E000000000000000000000000000;
                                 char22_4[36] <= 128'h0007E000000000000000000000000000;
                                 char22_4[37] <= 128'h0007E000000000000000000000000000;
                                 char22_4[38] <= 128'h0007E000000000000000000000000000;
                                 char22_4[39] <= 128'h0007E000000000000000000000000000;
                                 char22_4[40] <= 128'h0007E000000000000000000000000000;
                                 char22_4[41] <= 128'h0007E000000000000000000000000000;
                                 char22_4[42] <= 128'h0007E000000000000000000000000000;
                                 char22_4[43] <= 128'h0007E000000000000000000000000000;
                                 char22_4[44] <= 128'h0007E000000000000000000000000000;
                                 char22_4[45] <= 128'h0007E000000000000000000000000000;
                                 char22_4[46] <= 128'h0007E000000000000000000000000000;
                                 char22_4[47] <= 128'h0007E000000000000000000000000000;
                                 char22_4[48] <= 128'h0007E000000000000000000000000000;
                                 char22_4[49] <= 128'h0007E000000000000000000000000000;
                                 char22_4[50] <= 128'h0007E000000000000000000000000000;
                                 char22_4[51] <= 128'h000FF800000000000000000000000000;
                                 char22_4[52] <= 128'h03FFFFC0000000000000000000000000;
                                 char22_4[53] <= 128'h03FFFFC0000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//1
                           4'd2: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h001FFC00000000000000000000000000;
                                 char22_4[11] <= 128'h007FFF00000000000000000000000000;
                                 char22_4[12] <= 128'h01F83F80000000000000000000000000;
                                 char22_4[13] <= 128'h03E00FC0000000000000000000000000;
                                 char22_4[14] <= 128'h07C007E0000000000000000000000000;
                                 char22_4[15] <= 128'h078007E0000000000000000000000000;
                                 char22_4[16] <= 128'h0F8003F0000000000000000000000000;
                                 char22_4[17] <= 128'h0F8003F0000000000000000000000000;
                                 char22_4[18] <= 128'h1F8003F0000000000000000000000000;
                                 char22_4[19] <= 128'h1F8003F0000000000000000000000000;
                                 char22_4[20] <= 128'h1FC003F0000000000000000000000000;
                                 char22_4[21] <= 128'h1FC003F0000000000000000000000000;
                                 char22_4[22] <= 128'h1FC003F0000000000000000000000000;
                                 char22_4[23] <= 128'h0FC003F0000000000000000000000000;
                                 char22_4[24] <= 128'h07C003F0000000000000000000000000;
                                 char22_4[25] <= 128'h000003E0000000000000000000000000;
                                 char22_4[26] <= 128'h000007E0000000000000000000000000;
                                 char22_4[27] <= 128'h000007E0000000000000000000000000;
                                 char22_4[28] <= 128'h00000FC0000000000000000000000000;
                                 char22_4[29] <= 128'h00000F80000000000000000000000000;
                                 char22_4[30] <= 128'h00001F80000000000000000000000000;
                                 char22_4[31] <= 128'h00003F00000000000000000000000000;
                                 char22_4[32] <= 128'h00003E00000000000000000000000000;
                                 char22_4[33] <= 128'h00007C00000000000000000000000000;
                                 char22_4[34] <= 128'h0000F800000000000000000000000000;
                                 char22_4[35] <= 128'h0001F000000000000000000000000000;
                                 char22_4[36] <= 128'h0003E000000000000000000000000000;
                                 char22_4[37] <= 128'h0007C000000000000000000000000000;
                                 char22_4[38] <= 128'h000F8000000000000000000000000000;
                                 char22_4[39] <= 128'h001F0000000000000000000000000000;
                                 char22_4[40] <= 128'h003E0000000000000000000000000000;
                                 char22_4[41] <= 128'h007C0000000000000000000000000000;
                                 char22_4[42] <= 128'h00F80000000000000000000000000000;
                                 char22_4[43] <= 128'h01F00038000000000000000000000000;
                                 char22_4[44] <= 128'h01E00038000000000000000000000000;
                                 char22_4[45] <= 128'h03C00070000000000000000000000000;
                                 char22_4[46] <= 128'h07800070000000000000000000000000;
                                 char22_4[47] <= 128'h0F8000F0000000000000000000000000;
                                 char22_4[48] <= 128'h0F0000F0000000000000000000000000;
                                 char22_4[49] <= 128'h1E0003F0000000000000000000000000;
                                 char22_4[50] <= 128'h3FFFFFF0000000000000000000000000;
                                 char22_4[51] <= 128'h3FFFFFF0000000000000000000000000;
                                 char22_4[52] <= 128'h3FFFFFE0000000000000000000000000;
                                 char22_4[53] <= 128'h3FFFFFE0000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//2
                           4'd3: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h003FF000000000000000000000000000;
                                 char22_4[11] <= 128'h00FFFC00000000000000000000000000;
                                 char22_4[12] <= 128'h01F07E00000000000000000000000000;
                                 char22_4[13] <= 128'h03C03F00000000000000000000000000;
                                 char22_4[14] <= 128'h07801F80000000000000000000000000;
                                 char22_4[15] <= 128'h0F800FC0000000000000000000000000;
                                 char22_4[16] <= 128'h0F800FC0000000000000000000000000;
                                 char22_4[17] <= 128'h0F8007E0000000000000000000000000;
                                 char22_4[18] <= 128'h0FC007E0000000000000000000000000;
                                 char22_4[19] <= 128'h0FC007E0000000000000000000000000;
                                 char22_4[20] <= 128'h0FC007E0000000000000000000000000;
                                 char22_4[21] <= 128'h07C007E0000000000000000000000000;
                                 char22_4[22] <= 128'h000007E0000000000000000000000000;
                                 char22_4[23] <= 128'h000007E0000000000000000000000000;
                                 char22_4[24] <= 128'h000007C0000000000000000000000000;
                                 char22_4[25] <= 128'h00000FC0000000000000000000000000;
                                 char22_4[26] <= 128'h00000F80000000000000000000000000;
                                 char22_4[27] <= 128'h00001F00000000000000000000000000;
                                 char22_4[28] <= 128'h00007E00000000000000000000000000;
                                 char22_4[29] <= 128'h0003FC00000000000000000000000000;
                                 char22_4[30] <= 128'h001FF000000000000000000000000000;
                                 char22_4[31] <= 128'h001FFC00000000000000000000000000;
                                 char22_4[32] <= 128'h0000FF00000000000000000000000000;
                                 char22_4[33] <= 128'h00001F80000000000000000000000000;
                                 char22_4[34] <= 128'h00000FC0000000000000000000000000;
                                 char22_4[35] <= 128'h000007E0000000000000000000000000;
                                 char22_4[36] <= 128'h000003E0000000000000000000000000;
                                 char22_4[37] <= 128'h000003F0000000000000000000000000;
                                 char22_4[38] <= 128'h000003F0000000000000000000000000;
                                 char22_4[39] <= 128'h000001F0000000000000000000000000;
                                 char22_4[40] <= 128'h000001F8000000000000000000000000;
                                 char22_4[41] <= 128'h000001F8000000000000000000000000;
                                 char22_4[42] <= 128'h078001F8000000000000000000000000;
                                 char22_4[43] <= 128'h0FC001F8000000000000000000000000;
                                 char22_4[44] <= 128'h1FC001F8000000000000000000000000;
                                 char22_4[45] <= 128'h1FC003F0000000000000000000000000;
                                 char22_4[46] <= 128'h1FC003F0000000000000000000000000;
                                 char22_4[47] <= 128'h1FC003E0000000000000000000000000;
                                 char22_4[48] <= 128'h0F8007E0000000000000000000000000;
                                 char22_4[49] <= 128'h0F8007C0000000000000000000000000;
                                 char22_4[50] <= 128'h07C01F80000000000000000000000000;
                                 char22_4[51] <= 128'h03F07F00000000000000000000000000;
                                 char22_4[52] <= 128'h01FFFE00000000000000000000000000;
                                 char22_4[53] <= 128'h003FF000000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//3
                           4'd4: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h00001F00000000000000000000000000;
                                 char22_4[11] <= 128'h00001F00000000000000000000000000;
                                 char22_4[12] <= 128'h00003F00000000000000000000000000;
                                 char22_4[13] <= 128'h00003F00000000000000000000000000;
                                 char22_4[14] <= 128'h00007F00000000000000000000000000;
                                 char22_4[15] <= 128'h0000FF00000000000000000000000000;
                                 char22_4[16] <= 128'h0000FF00000000000000000000000000;
                                 char22_4[17] <= 128'h0001FF00000000000000000000000000;
                                 char22_4[18] <= 128'h0003FF00000000000000000000000000;
                                 char22_4[19] <= 128'h0003BF00000000000000000000000000;
                                 char22_4[20] <= 128'h0007BF00000000000000000000000000;
                                 char22_4[21] <= 128'h00073F00000000000000000000000000;
                                 char22_4[22] <= 128'h000F3F00000000000000000000000000;
                                 char22_4[23] <= 128'h001E3F00000000000000000000000000;
                                 char22_4[24] <= 128'h001C3F00000000000000000000000000;
                                 char22_4[25] <= 128'h003C3F00000000000000000000000000;
                                 char22_4[26] <= 128'h00783F00000000000000000000000000;
                                 char22_4[27] <= 128'h00783F00000000000000000000000000;
                                 char22_4[28] <= 128'h00F03F00000000000000000000000000;
                                 char22_4[29] <= 128'h00E03F00000000000000000000000000;
                                 char22_4[30] <= 128'h01E03F00000000000000000000000000;
                                 char22_4[31] <= 128'h03C03F00000000000000000000000000;
                                 char22_4[32] <= 128'h03803F00000000000000000000000000;
                                 char22_4[33] <= 128'h07803F00000000000000000000000000;
                                 char22_4[34] <= 128'h0F003F00000000000000000000000000;
                                 char22_4[35] <= 128'h0F003F00000000000000000000000000;
                                 char22_4[36] <= 128'h1E003F00000000000000000000000000;
                                 char22_4[37] <= 128'h1C003F00000000000000000000000000;
                                 char22_4[38] <= 128'h3C003F00000000000000000000000000;
                                 char22_4[39] <= 128'h7FFFFFFE000000000000000000000000;
                                 char22_4[40] <= 128'h7FFFFFFE000000000000000000000000;
                                 char22_4[41] <= 128'h00003F00000000000000000000000000;
                                 char22_4[42] <= 128'h00003F00000000000000000000000000;
                                 char22_4[43] <= 128'h00003F00000000000000000000000000;
                                 char22_4[44] <= 128'h00003F00000000000000000000000000;
                                 char22_4[45] <= 128'h00003F00000000000000000000000000;
                                 char22_4[46] <= 128'h00003F00000000000000000000000000;
                                 char22_4[47] <= 128'h00003F00000000000000000000000000;
                                 char22_4[48] <= 128'h00003F00000000000000000000000000;
                                 char22_4[49] <= 128'h00003F00000000000000000000000000;
                                 char22_4[50] <= 128'h00003F00000000000000000000000000;
                                 char22_4[51] <= 128'h00007F80000000000000000000000000;
                                 char22_4[52] <= 128'h000FFFFC000000000000000000000000;
                                 char22_4[53] <= 128'h000FFFFC000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//4
                           4'd5: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h00000000000000000000000000000000;
                                 char22_4[11] <= 128'h03FFFFF0000000000000000000000000;
                                 char22_4[12] <= 128'h03FFFFF0000000000000000000000000;
                                 char22_4[13] <= 128'h03FFFFF0000000000000000000000000;
                                 char22_4[14] <= 128'h03FFFFE0000000000000000000000000;
                                 char22_4[15] <= 128'h03800000000000000000000000000000;
                                 char22_4[16] <= 128'h03800000000000000000000000000000;
                                 char22_4[17] <= 128'h03800000000000000000000000000000;
                                 char22_4[18] <= 128'h03800000000000000000000000000000;
                                 char22_4[19] <= 128'h03800000000000000000000000000000;
                                 char22_4[20] <= 128'h07800000000000000000000000000000;
                                 char22_4[21] <= 128'h07800000000000000000000000000000;
                                 char22_4[22] <= 128'h07800000000000000000000000000000;
                                 char22_4[23] <= 128'h07800000000000000000000000000000;
                                 char22_4[24] <= 128'h07800000000000000000000000000000;
                                 char22_4[25] <= 128'h07800000000000000000000000000000;
                                 char22_4[26] <= 128'h078FF800000000000000000000000000;
                                 char22_4[27] <= 128'h073FFE00000000000000000000000000;
                                 char22_4[28] <= 128'h077FFF80000000000000000000000000;
                                 char22_4[29] <= 128'h07FC3F80000000000000000000000000;
                                 char22_4[30] <= 128'h07E00FC0000000000000000000000000;
                                 char22_4[31] <= 128'h07C007E0000000000000000000000000;
                                 char22_4[32] <= 128'h078007E0000000000000000000000000;
                                 char22_4[33] <= 128'h078003F0000000000000000000000000;
                                 char22_4[34] <= 128'h000003F0000000000000000000000000;
                                 char22_4[35] <= 128'h000001F0000000000000000000000000;
                                 char22_4[36] <= 128'h000001F8000000000000000000000000;
                                 char22_4[37] <= 128'h000001F8000000000000000000000000;
                                 char22_4[38] <= 128'h000001F8000000000000000000000000;
                                 char22_4[39] <= 128'h000001F8000000000000000000000000;
                                 char22_4[40] <= 128'h000001F8000000000000000000000000;
                                 char22_4[41] <= 128'h078001F8000000000000000000000000;
                                 char22_4[42] <= 128'h0FC001F8000000000000000000000000;
                                 char22_4[43] <= 128'h1FC001F0000000000000000000000000;
                                 char22_4[44] <= 128'h1FC001F0000000000000000000000000;
                                 char22_4[45] <= 128'h1FC003F0000000000000000000000000;
                                 char22_4[46] <= 128'h1F8003F0000000000000000000000000;
                                 char22_4[47] <= 128'h1F8003E0000000000000000000000000;
                                 char22_4[48] <= 128'h0F8007E0000000000000000000000000;
                                 char22_4[49] <= 128'h078007C0000000000000000000000000;
                                 char22_4[50] <= 128'h07C01F80000000000000000000000000;
                                 char22_4[51] <= 128'h03F83F00000000000000000000000000;
                                 char22_4[52] <= 128'h00FFFE00000000000000000000000000;
                                 char22_4[53] <= 128'h003FF800000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//5
                           4'd6: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h0007FE00000000000000000000000000;
                                 char22_4[11] <= 128'h001FFF80000000000000000000000000;
                                 char22_4[12] <= 128'h003F0FC0000000000000000000000000;
                                 char22_4[13] <= 128'h007C07C0000000000000000000000000;
                                 char22_4[14] <= 128'h00F807E0000000000000000000000000;
                                 char22_4[15] <= 128'h01F007E0000000000000000000000000;
                                 char22_4[16] <= 128'h03E007E0000000000000000000000000;
                                 char22_4[17] <= 128'h03C007E0000000000000000000000000;
                                 char22_4[18] <= 128'h07C003C0000000000000000000000000;
                                 char22_4[19] <= 128'h07C00000000000000000000000000000;
                                 char22_4[20] <= 128'h0FC00000000000000000000000000000;
                                 char22_4[21] <= 128'h0F800000000000000000000000000000;
                                 char22_4[22] <= 128'h0F800000000000000000000000000000;
                                 char22_4[23] <= 128'h1F800000000000000000000000000000;
                                 char22_4[24] <= 128'h1F800000000000000000000000000000;
                                 char22_4[25] <= 128'h1F800000000000000000000000000000;
                                 char22_4[26] <= 128'h1F87FE00000000000000000000000000;
                                 char22_4[27] <= 128'h1F9FFF80000000000000000000000000;
                                 char22_4[28] <= 128'h1FBFFFC0000000000000000000000000;
                                 char22_4[29] <= 128'h3FFE1FC0000000000000000000000000;
                                 char22_4[30] <= 128'h3FF807E0000000000000000000000000;
                                 char22_4[31] <= 128'h3FE003F0000000000000000000000000;
                                 char22_4[32] <= 128'h3FE003F0000000000000000000000000;
                                 char22_4[33] <= 128'h3FC001F8000000000000000000000000;
                                 char22_4[34] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[35] <= 128'h3F8001F8000000000000000000000000;
                                 char22_4[36] <= 128'h3F8000F8000000000000000000000000;
                                 char22_4[37] <= 128'h3F8000F8000000000000000000000000;
                                 char22_4[38] <= 128'h3F8000F8000000000000000000000000;
                                 char22_4[39] <= 128'h1F8000F8000000000000000000000000;
                                 char22_4[40] <= 128'h1F8000F8000000000000000000000000;
                                 char22_4[41] <= 128'h1F8000F8000000000000000000000000;
                                 char22_4[42] <= 128'h1F8000F8000000000000000000000000;
                                 char22_4[43] <= 128'h1F8000F8000000000000000000000000;
                                 char22_4[44] <= 128'h0FC001F8000000000000000000000000;
                                 char22_4[45] <= 128'h0FC001F8000000000000000000000000;
                                 char22_4[46] <= 128'h0FC001F0000000000000000000000000;
                                 char22_4[47] <= 128'h07E001F0000000000000000000000000;
                                 char22_4[48] <= 128'h03E003E0000000000000000000000000;
                                 char22_4[49] <= 128'h03F003E0000000000000000000000000;
                                 char22_4[50] <= 128'h01F807C0000000000000000000000000;
                                 char22_4[51] <= 128'h00FE1F80000000000000000000000000;
                                 char22_4[52] <= 128'h007FFE00000000000000000000000000;
                                 char22_4[53] <= 128'h001FF800000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//6
                           4'd7: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h00000000000000000000000000000000;
                                 char22_4[11] <= 128'h07FFFFF8000000000000000000000000;
                                 char22_4[12] <= 128'h07FFFFF8000000000000000000000000;
                                 char22_4[13] <= 128'h07FFFFF8000000000000000000000000;
                                 char22_4[14] <= 128'h0FFFFFF0000000000000000000000000;
                                 char22_4[15] <= 128'h0FC000E0000000000000000000000000;
                                 char22_4[16] <= 128'h0F8001E0000000000000000000000000;
                                 char22_4[17] <= 128'h0F0001C0000000000000000000000000;
                                 char22_4[18] <= 128'h0E0003C0000000000000000000000000;
                                 char22_4[19] <= 128'h0E000780000000000000000000000000;
                                 char22_4[20] <= 128'h1E000780000000000000000000000000;
                                 char22_4[21] <= 128'h1C000F00000000000000000000000000;
                                 char22_4[22] <= 128'h00000F00000000000000000000000000;
                                 char22_4[23] <= 128'h00001E00000000000000000000000000;
                                 char22_4[24] <= 128'h00001E00000000000000000000000000;
                                 char22_4[25] <= 128'h00003C00000000000000000000000000;
                                 char22_4[26] <= 128'h00003C00000000000000000000000000;
                                 char22_4[27] <= 128'h00007800000000000000000000000000;
                                 char22_4[28] <= 128'h00007800000000000000000000000000;
                                 char22_4[29] <= 128'h0000F800000000000000000000000000;
                                 char22_4[30] <= 128'h0000F000000000000000000000000000;
                                 char22_4[31] <= 128'h0001F000000000000000000000000000;
                                 char22_4[32] <= 128'h0001E000000000000000000000000000;
                                 char22_4[33] <= 128'h0003E000000000000000000000000000;
                                 char22_4[34] <= 128'h0003E000000000000000000000000000;
                                 char22_4[35] <= 128'h0003E000000000000000000000000000;
                                 char22_4[36] <= 128'h0007C000000000000000000000000000;
                                 char22_4[37] <= 128'h0007C000000000000000000000000000;
                                 char22_4[38] <= 128'h0007C000000000000000000000000000;
                                 char22_4[39] <= 128'h000FC000000000000000000000000000;
                                 char22_4[40] <= 128'h000FC000000000000000000000000000;
                                 char22_4[41] <= 128'h000FC000000000000000000000000000;
                                 char22_4[42] <= 128'h000FC000000000000000000000000000;
                                 char22_4[43] <= 128'h001FC000000000000000000000000000;
                                 char22_4[44] <= 128'h001FC000000000000000000000000000;
                                 char22_4[45] <= 128'h001FC000000000000000000000000000;
                                 char22_4[46] <= 128'h001FC000000000000000000000000000;
                                 char22_4[47] <= 128'h001FC000000000000000000000000000;
                                 char22_4[48] <= 128'h001FC000000000000000000000000000;
                                 char22_4[49] <= 128'h001FC000000000000000000000000000;
                                 char22_4[50] <= 128'h001FC000000000000000000000000000;
                                 char22_4[51] <= 128'h001FC000000000000000000000000000;
                                 char22_4[52] <= 128'h001FC000000000000000000000000000;
                                 char22_4[53] <= 128'h000F8000000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//7
                           4'd8: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h003FF800000000000000000000000000;
                                 char22_4[11] <= 128'h00FFFE00000000000000000000000000;
                                 char22_4[12] <= 128'h01F81F80000000000000000000000000;
                                 char22_4[13] <= 128'h03E00FC0000000000000000000000000;
                                 char22_4[14] <= 128'h07C003E0000000000000000000000000;
                                 char22_4[15] <= 128'h0F8003E0000000000000000000000000;
                                 char22_4[16] <= 128'h0F8001F0000000000000000000000000;
                                 char22_4[17] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[18] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[19] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[20] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[21] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[22] <= 128'h1F8001F0000000000000000000000000;
                                 char22_4[23] <= 128'h1FC001F0000000000000000000000000;
                                 char22_4[24] <= 128'h0FC001F0000000000000000000000000;
                                 char22_4[25] <= 128'h0FF003E0000000000000000000000000;
                                 char22_4[26] <= 128'h07F803C0000000000000000000000000;
                                 char22_4[27] <= 128'h03FE0F80000000000000000000000000;
                                 char22_4[28] <= 128'h01FF9F00000000000000000000000000;
                                 char22_4[29] <= 128'h00FFFE00000000000000000000000000;
                                 char22_4[30] <= 128'h003FF800000000000000000000000000;
                                 char22_4[31] <= 128'h007FFC00000000000000000000000000;
                                 char22_4[32] <= 128'h01F7FF00000000000000000000000000;
                                 char22_4[33] <= 128'h03E1FF80000000000000000000000000;
                                 char22_4[34] <= 128'h07C07FC0000000000000000000000000;
                                 char22_4[35] <= 128'h0F801FE0000000000000000000000000;
                                 char22_4[36] <= 128'h0F800FE0000000000000000000000000;
                                 char22_4[37] <= 128'h1F0007F0000000000000000000000000;
                                 char22_4[38] <= 128'h1F0003F0000000000000000000000000;
                                 char22_4[39] <= 128'h3E0001F8000000000000000000000000;
                                 char22_4[40] <= 128'h3E0001F8000000000000000000000000;
                                 char22_4[41] <= 128'h3E0001F8000000000000000000000000;
                                 char22_4[42] <= 128'h3E0000F8000000000000000000000000;
                                 char22_4[43] <= 128'h3E0000F8000000000000000000000000;
                                 char22_4[44] <= 128'h3E0000F8000000000000000000000000;
                                 char22_4[45] <= 128'h3E0000F8000000000000000000000000;
                                 char22_4[46] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[47] <= 128'h1F0001F0000000000000000000000000;
                                 char22_4[48] <= 128'h0F8003E0000000000000000000000000;
                                 char22_4[49] <= 128'h0FC003E0000000000000000000000000;
                                 char22_4[50] <= 128'h07E007C0000000000000000000000000;
                                 char22_4[51] <= 128'h01F83F80000000000000000000000000;
                                 char22_4[52] <= 128'h00FFFE00000000000000000000000000;
                                 char22_4[53] <= 128'h003FF800000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//8
                           4'd9: begin
                                 char22_4[0] <= 128'h00000000000000000000000000000000;
                                 char22_4[1] <= 128'h00000000000000000000000000000000;
                                 char22_4[2] <= 128'h00000000000000000000000000000000;
                                 char22_4[3] <= 128'h00000000000000000000000000000000;
                                 char22_4[4] <= 128'h00000000000000000000000000000000;
                                 char22_4[5] <= 128'h00000000000000000000000000000000;
                                 char22_4[6] <= 128'h00000000000000000000000000000000;
                                 char22_4[7] <= 128'h00000000000000000000000000000000;
                                 char22_4[8] <= 128'h00000000000000000000000000000000;
                                 char22_4[9] <= 128'h00000000000000000000000000000000;
                                 char22_4[10] <= 128'h003FF000000000000000000000000000;
                                 char22_4[11] <= 128'h00FFFC00000000000000000000000000;
                                 char22_4[12] <= 128'h01F83F00000000000000000000000000;
                                 char22_4[13] <= 128'h03E01F80000000000000000000000000;
                                 char22_4[14] <= 128'h07C00F80000000000000000000000000;
                                 char22_4[15] <= 128'h0FC007C0000000000000000000000000;
                                 char22_4[16] <= 128'h0F8003E0000000000000000000000000;
                                 char22_4[17] <= 128'h1F8003E0000000000000000000000000;
                                 char22_4[18] <= 128'h1F0003F0000000000000000000000000;
                                 char22_4[19] <= 128'h1F0003F0000000000000000000000000;
                                 char22_4[20] <= 128'h3F0001F0000000000000000000000000;
                                 char22_4[21] <= 128'h3F0001F0000000000000000000000000;
                                 char22_4[22] <= 128'h3F0001F8000000000000000000000000;
                                 char22_4[23] <= 128'h3F0001F8000000000000000000000000;
                                 char22_4[24] <= 128'h3F0001F8000000000000000000000000;
                                 char22_4[25] <= 128'h3F0001F8000000000000000000000000;
                                 char22_4[26] <= 128'h3F0001F8000000000000000000000000;
                                 char22_4[27] <= 128'h3F0001F8000000000000000000000000;
                                 char22_4[28] <= 128'h3F0003F8000000000000000000000000;
                                 char22_4[29] <= 128'h1F8003F8000000000000000000000000;
                                 char22_4[30] <= 128'h1F8007F8000000000000000000000000;
                                 char22_4[31] <= 128'h1F800FF8000000000000000000000000;
                                 char22_4[32] <= 128'h0FC01FF8000000000000000000000000;
                                 char22_4[33] <= 128'h0FE03FF8000000000000000000000000;
                                 char22_4[34] <= 128'h07F8FDF8000000000000000000000000;
                                 char22_4[35] <= 128'h03FFF9F8000000000000000000000000;
                                 char22_4[36] <= 128'h01FFF1F8000000000000000000000000;
                                 char22_4[37] <= 128'h003F83F8000000000000000000000000;
                                 char22_4[38] <= 128'h000003F0000000000000000000000000;
                                 char22_4[39] <= 128'h000003F0000000000000000000000000;
                                 char22_4[40] <= 128'h000003F0000000000000000000000000;
                                 char22_4[41] <= 128'h000003F0000000000000000000000000;
                                 char22_4[42] <= 128'h000007E0000000000000000000000000;
                                 char22_4[43] <= 128'h000007E0000000000000000000000000;
                                 char22_4[44] <= 128'h000007C0000000000000000000000000;
                                 char22_4[45] <= 128'h03C007C0000000000000000000000000;
                                 char22_4[46] <= 128'h07C00F80000000000000000000000000;
                                 char22_4[47] <= 128'h0FE00F80000000000000000000000000;
                                 char22_4[48] <= 128'h0FE01F00000000000000000000000000;
                                 char22_4[49] <= 128'h0FE03E00000000000000000000000000;
                                 char22_4[50] <= 128'h07E07E00000000000000000000000000;
                                 char22_4[51] <= 128'h07F1F800000000000000000000000000;
                                 char22_4[52] <= 128'h03FFF000000000000000000000000000;
                                 char22_4[53] <= 128'h00FFC000000000000000000000000000;
                                 char22_4[54] <= 128'h00000000000000000000000000000000;
                                 char22_4[55] <= 128'h00000000000000000000000000000000;
                                 char22_4[56] <= 128'h00000000000000000000000000000000;
                                 char22_4[57] <= 128'h00000000000000000000000000000000;
                                 char22_4[58] <= 128'h00000000000000000000000000000000;
                                 char22_4[59] <= 128'h00000000000000000000000000000000;
                                 char22_4[60] <= 128'h00000000000000000000000000000000;
                                 char22_4[61] <= 128'h00000000000000000000000000000000;
                                 char22_4[62] <= 128'h00000000000000000000000000000000;
                                 char22_4[63] <= 128'h00000000000000000000000000000000;
                           end//9
                           default: begin
                               char22_4[0] <= char22_4[0];
                               char22_4[1] <= char22_4[1];
                               char22_4[2] <= char22_4[2];
                               char22_4[3] <= char22_4[3];
                               char22_4[4] <= char22_4[4];
                               char22_4[5] <= char22_4[5];
                               char22_4[6] <= char22_4[6];
                               char22_4[7] <= char22_4[7];
                               char22_4[8] <= char22_4[8];
                               char22_4[9] <= char22_4[9];
                               char22_4[10] <= char22_4[10];
                               char22_4[11] <= char22_4[11];
                               char22_4[12] <= char22_4[12];
                               char22_4[13] <= char22_4[13];
                               char22_4[14] <= char22_4[14];
                               char22_4[15] <= char22_4[15];
                               char22_4[16] <= char22_4[16];
                               char22_4[17] <= char22_4[17];
                               char22_4[18] <= char22_4[18];
                               char22_4[19] <= char22_4[19];
                               char22_4[20] <= char22_4[20];
                               char22_4[21] <= char22_4[21];
                               char22_4[22] <= char22_4[22];
                               char22_4[23] <= char22_4[23];
                               char22_4[24] <= char22_4[24];
                               char22_4[25] <= char22_4[25];
                               char22_4[26] <= char22_4[26];
                               char22_4[27] <= char22_4[27];
                               char22_4[28] <= char22_4[28];
                               char22_4[29] <= char22_4[29];
                               char22_4[30] <= char22_4[30];
                               char22_4[31] <= char22_4[31];
                               char22_4[32] <= char22_4[32];
                               char22_4[33] <= char22_4[33];
                               char22_4[34] <= char22_4[34];
                               char22_4[35] <= char22_4[35];
                               char22_4[36] <= char22_4[36];
                               char22_4[37] <= char22_4[37];
                               char22_4[38] <= char22_4[38];
                               char22_4[39] <= char22_4[39];
                               char22_4[40] <= char22_4[40];
                               char22_4[41] <= char22_4[41];
                               char22_4[42] <= char22_4[42];
                               char22_4[43] <= char22_4[43];
                               char22_4[44] <= char22_4[44];
                               char22_4[45] <= char22_4[45];
                               char22_4[46] <= char22_4[46];
                               char22_4[47] <= char22_4[47];
                               char22_4[48] <= char22_4[48];
                               char22_4[49] <= char22_4[49];
                               char22_4[50] <= char22_4[50];
                               char22_4[51] <= char22_4[51];
                               char22_4[52] <= char22_4[52];
                               char22_4[53] <= char22_4[53];
                               char22_4[54] <= char22_4[54];
                               char22_4[55] <= char22_4[55];
                               char22_4[56] <= char22_4[56];
                               char22_4[57] <= char22_4[57];
                               char22_4[58] <= char22_4[58];
                               char22_4[59] <= char22_4[59];
                               char22_4[60] <= char22_4[60];
                               char22_4[61] <= char22_4[61];
                               char22_4[62] <= char22_4[62];
                               char22_4[63] <= char22_4[63];
                           end
                       endcase
               
         case(a1/w1)
                           4'd0: begin
                               char33_0[  0] <= 32'h00000000;
                               char33_0[  1] <= 32'h00000000;
                               char33_0[  2] <= 32'h00000000;
                               char33_0[  3] <= 32'h00000000;
                               char33_0[  4] <= 32'h00000000;
                               char33_0[  5] <= 32'h00000000;
                               char33_0[  6] <= 32'h00000000;
                               char33_0[  7] <= 32'h00000000;
                               char33_0[  8] <= 32'h00000000;
                               char33_0[  9] <= 32'h00000000;
                               char33_0[10] <= 32'h000FF000;
                               char33_0[11] <= 32'h003FFC00;
                               char33_0[12] <= 32'h007E7E00;
                               char33_0[13] <= 32'h00F81F00;
                               char33_0[14] <= 32'h01F00F80;
                               char33_0[15] <= 32'h03F00FC0;
                               char33_0[16] <= 32'h03E007C0;
                               char33_0[17] <= 32'h07E007E0;
                               char33_0[18] <= 32'h07C003E0;
                               char33_0[19] <= 32'h0FC003F0;
                               char33_0[20] <= 32'h0FC003F0;
                               char33_0[21] <= 32'h0FC003F0;
                               char33_0[22] <= 32'h1F8001F8;
                               char33_0[23] <= 32'h1F8001F8;
                               char33_0[24] <= 32'h1F8001F8;
                               char33_0[25] <= 32'h1F8001F8;
                               char33_0[26] <= 32'h1F8001F8;
                               char33_0[27] <= 32'h3F8001F8;
                               char33_0[28] <= 32'h3F8001F8;
                               char33_0[29] <= 32'h3F8001F8;
                               char33_0[30] <= 32'h3F8001F8;
                               char33_0[31] <= 32'h3F8001F8;
                               char33_0[32] <= 32'h3F8001F8;
                               char33_0[33] <= 32'h3F8001F8;
                               char33_0[34] <= 32'h3F8001F8;
                               char33_0[35] <= 32'h3F8001F8;
                               char33_0[36] <= 32'h3F8001F8;
                               char33_0[37] <= 32'h1F8001F8;
                               char33_0[38] <= 32'h1F8001F8;
                               char33_0[39] <= 32'h1F8001F8;
                               char33_0[40] <= 32'h1F8001F8;
                               char33_0[41] <= 32'h1F8001F0;
                               char33_0[42] <= 32'h0F8003F0;
                               char33_0[43] <= 32'h0FC003F0;
                               char33_0[44] <= 32'h0FC003F0;
                               char33_0[45] <= 32'h07C003E0;
                               char33_0[46] <= 32'h07E007E0;
                               char33_0[47] <= 32'h03E007C0;
                               char33_0[48] <= 32'h03F00FC0;
                               char33_0[49] <= 32'h01F00F80;
                               char33_0[50] <= 32'h00F81F00;
                               char33_0[51] <= 32'h007E7E00;
                               char33_0[52] <= 32'h003FFC00;
                               char33_0[53] <= 32'h000FF000;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//0
                           4'd1: begin
                               char33_0[  0] <= 32'h00000000;
                               char33_0[  1] <= 32'h00000000;
                               char33_0[  2] <= 32'h00000000;
                               char33_0[  3] <= 32'h00000000;
                               char33_0[  4] <= 32'h00000000;
                               char33_0[  5] <= 32'h00000000;
                               char33_0[  6] <= 32'h00000000;
                               char33_0[  7] <= 32'h00000000;
                               char33_0[  8] <= 32'h00000000;
                               char33_0[  9] <= 32'h00000000;
                               char33_0[10] <= 32'h0000E000;
                               char33_0[11] <= 32'h0001E000;
                               char33_0[12] <= 32'h0003E000;
                               char33_0[13] <= 32'h001FE000;
                               char33_0[14] <= 32'h03FFE000;
                               char33_0[15] <= 32'h03FFE000;
                               char33_0[16] <= 32'h0007E000;
                               char33_0[17] <= 32'h0007E000;
                               char33_0[18] <= 32'h0007E000;
                               char33_0[19] <= 32'h0007E000;
                               char33_0[20] <= 32'h0007E000;
                               char33_0[21] <= 32'h0007E000;
                               char33_0[22] <= 32'h0007E000;
                               char33_0[23] <= 32'h0007E000;
                               char33_0[24] <= 32'h0007E000;
                               char33_0[25] <= 32'h0007E000;
                               char33_0[26] <= 32'h0007E000;
                               char33_0[27] <= 32'h0007E000;
                               char33_0[28] <= 32'h0007E000;
                               char33_0[29] <= 32'h0007E000;
                               char33_0[30] <= 32'h0007E000;
                               char33_0[31] <= 32'h0007E000;
                               char33_0[32] <= 32'h0007E000;
                               char33_0[33] <= 32'h0007E000;
                               char33_0[34] <= 32'h0007E000;
                               char33_0[35] <= 32'h0007E000;
                               char33_0[36] <= 32'h0007E000;
                               char33_0[37] <= 32'h0007E000;
                               char33_0[38] <= 32'h0007E000;
                               char33_0[39] <= 32'h0007E000;
                               char33_0[40] <= 32'h0007E000;
                               char33_0[41] <= 32'h0007E000;
                               char33_0[42] <= 32'h0007E000;
                               char33_0[43] <= 32'h0007E000;
                               char33_0[44] <= 32'h0007E000;
                               char33_0[45] <= 32'h0007E000;
                               char33_0[46] <= 32'h0007E000;
                               char33_0[47] <= 32'h0007E000;
                               char33_0[48] <= 32'h0007E000;
                               char33_0[49] <= 32'h0007E000;
                               char33_0[50] <= 32'h0007E000;
                               char33_0[51] <= 32'h000FF800;
                               char33_0[52] <= 32'h03FFFFC0;
                               char33_0[53] <= 32'h03FFFFC0;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//1
                           4'd2: begin
                               char33_0[  0] <= 32'h00000000;
                               char33_0[  1] <= 32'h00000000;
                               char33_0[  2] <= 32'h00000000;
                               char33_0[  3] <= 32'h00000000;
                               char33_0[  4] <= 32'h00000000;
                               char33_0[  5] <= 32'h00000000;
                               char33_0[  6] <= 32'h00000000;
                               char33_0[  7] <= 32'h00000000;
                               char33_0[  8] <= 32'h00000000;
                               char33_0[  9] <= 32'h00000000;
                               char33_0[10] <= 32'h001FFC00;
                               char33_0[11] <= 32'h007FFF00;
                               char33_0[12] <= 32'h01F83F80;
                               char33_0[13] <= 32'h03E00FC0;
                               char33_0[14] <= 32'h07C007E0;
                               char33_0[15] <= 32'h078007E0;
                               char33_0[16] <= 32'h0F8003F0;
                               char33_0[17] <= 32'h0F8003F0;
                               char33_0[18] <= 32'h1F8003F0;
                               char33_0[19] <= 32'h1F8003F0;
                               char33_0[20] <= 32'h1FC003F0;
                               char33_0[21] <= 32'h1FC003F0;
                               char33_0[22] <= 32'h1FC003F0;
                               char33_0[23] <= 32'h0FC003F0;
                               char33_0[24] <= 32'h07C003F0;
                               char33_0[25] <= 32'h000003E0;
                               char33_0[26] <= 32'h000007E0;
                               char33_0[27] <= 32'h000007E0;
                               char33_0[28] <= 32'h00000FC0;
                               char33_0[29] <= 32'h00000F80;
                               char33_0[30] <= 32'h00001F80;
                               char33_0[31] <= 32'h00003F00;
                               char33_0[32] <= 32'h00003E00;
                               char33_0[33] <= 32'h00007C00;
                               char33_0[34] <= 32'h0000F800;
                               char33_0[35] <= 32'h0001F000;
                               char33_0[36] <= 32'h0003E000;
                               char33_0[37] <= 32'h0007C000;
                               char33_0[38] <= 32'h000F8000;
                               char33_0[39] <= 32'h001F0000;
                               char33_0[40] <= 32'h003E0000;
                               char33_0[41] <= 32'h007C0000;
                               char33_0[42] <= 32'h00F80000;
                               char33_0[43] <= 32'h01F00038;
                               char33_0[44] <= 32'h01E00038;
                               char33_0[45] <= 32'h03C00070;
                               char33_0[46] <= 32'h07800070;
                               char33_0[47] <= 32'h0F8000F0;
                               char33_0[48] <= 32'h0F0000F0;
                               char33_0[49] <= 32'h1E0003F0;
                               char33_0[50] <= 32'h3FFFFFF0;
                               char33_0[51] <= 32'h3FFFFFF0;
                               char33_0[52] <= 32'h3FFFFFE0;
                               char33_0[53] <= 32'h3FFFFFE0;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//2
                           4'd3: begin
                               char33_0[  0] <= 32'h00000000;
                               char33_0[  1] <= 32'h00000000;
                               char33_0[  2] <= 32'h00000000;
                               char33_0[  3] <= 32'h00000000;
                               char33_0[  4] <= 32'h00000000;
                               char33_0[  5] <= 32'h00000000;
                               char33_0[  6] <= 32'h00000000;
                               char33_0[  7] <= 32'h00000000;
                               char33_0[  8] <= 32'h00000000;
                               char33_0[  9] <= 32'h00000000;
                               char33_0[10] <= 32'h003FF000;
                               char33_0[11] <= 32'h00FFFC00;
                               char33_0[12] <= 32'h01F07E00;
                               char33_0[13] <= 32'h03C03F00;
                               char33_0[14] <= 32'h07801F80;
                               char33_0[15] <= 32'h0F800FC0;
                               char33_0[16] <= 32'h0F800FC0;
                               char33_0[17] <= 32'h0F8007E0;
                               char33_0[18] <= 32'h0FC007E0;
                               char33_0[19] <= 32'h0FC007E0;
                               char33_0[20] <= 32'h0FC007E0;
                               char33_0[21] <= 32'h07C007E0;
                               char33_0[22] <= 32'h000007E0;
                               char33_0[23] <= 32'h000007E0;
                               char33_0[24] <= 32'h000007C0;
                               char33_0[25] <= 32'h00000FC0;
                               char33_0[26] <= 32'h00000F80;
                               char33_0[27] <= 32'h00001F00;
                               char33_0[28] <= 32'h00007E00;
                               char33_0[29] <= 32'h0003FC00;
                               char33_0[30] <= 32'h001FF000;
                               char33_0[31] <= 32'h001FFC00;
                               char33_0[32] <= 32'h0000FF00;
                               char33_0[33] <= 32'h00001F80;
                               char33_0[34] <= 32'h00000FC0;
                               char33_0[35] <= 32'h000007E0;
                               char33_0[36] <= 32'h000003E0;
                               char33_0[37] <= 32'h000003F0;
                               char33_0[38] <= 32'h000003F0;
                               char33_0[39] <= 32'h000001F0;
                               char33_0[40] <= 32'h000001F8;
                               char33_0[41] <= 32'h000001F8;
                               char33_0[42] <= 32'h078001F8;
                               char33_0[43] <= 32'h0FC001F8;
                               char33_0[44] <= 32'h1FC001F8;
                               char33_0[45] <= 32'h1FC003F0;
                               char33_0[46] <= 32'h1FC003F0;
                               char33_0[47] <= 32'h1FC003E0;
                               char33_0[48] <= 32'h0F8007E0;
                               char33_0[49] <= 32'h0F8007C0;
                               char33_0[50] <= 32'h07C01F80;
                               char33_0[51] <= 32'h03F07F00;
                               char33_0[52] <= 32'h01FFFE00;
                               char33_0[53] <= 32'h003FF000;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//3
                           4'd4: begin
                               char33_0[  0] <= 32'h00000000;
                               char33_0[  1] <= 32'h00000000;
                               char33_0[  2] <= 32'h00000000;
                               char33_0[  3] <= 32'h00000000;
                               char33_0[  4] <= 32'h00000000;
                               char33_0[  5] <= 32'h00000000;
                               char33_0[  6] <= 32'h00000000;
                               char33_0[  7] <= 32'h00000000;
                               char33_0[  8] <= 32'h00000000;
                               char33_0[  9] <= 32'h00000000;
                               char33_0[10] <= 32'h00001F00;
                               char33_0[11] <= 32'h00001F00;
                               char33_0[12] <= 32'h00003F00;
                               char33_0[13] <= 32'h00003F00;
                               char33_0[14] <= 32'h00007F00;
                               char33_0[15] <= 32'h0000FF00;
                               char33_0[16] <= 32'h0000FF00;
                               char33_0[17] <= 32'h0001FF00;
                               char33_0[18] <= 32'h0003FF00;
                               char33_0[19] <= 32'h0003BF00;
                               char33_0[20] <= 32'h0007BF00;
                               char33_0[21] <= 32'h00073F00;
                               char33_0[22] <= 32'h000F3F00;
                               char33_0[23] <= 32'h001E3F00;
                               char33_0[24] <= 32'h001C3F00;
                               char33_0[25] <= 32'h003C3F00;
                               char33_0[26] <= 32'h00783F00;
                               char33_0[27] <= 32'h00783F00;
                               char33_0[28] <= 32'h00F03F00;
                               char33_0[29] <= 32'h00E03F00;
                               char33_0[30] <= 32'h01E03F00;
                               char33_0[31] <= 32'h03C03F00;
                               char33_0[32] <= 32'h03803F00;
                               char33_0[33] <= 32'h07803F00;
                               char33_0[34] <= 32'h0F003F00;
                               char33_0[35] <= 32'h0F003F00;
                               char33_0[36] <= 32'h1E003F00;
                               char33_0[37] <= 32'h1C003F00;
                               char33_0[38] <= 32'h3C003F00;
                               char33_0[39] <= 32'h7FFFFFFE;
                               char33_0[40] <= 32'h7FFFFFFE;
                               char33_0[41] <= 32'h00003F00;
                               char33_0[42] <= 32'h00003F00;
                               char33_0[43] <= 32'h00003F00;
                               char33_0[44] <= 32'h00003F00;
                               char33_0[45] <= 32'h00003F00;
                               char33_0[46] <= 32'h00003F00;
                               char33_0[47] <= 32'h00003F00;
                               char33_0[48] <= 32'h00003F00;
                               char33_0[49] <= 32'h00003F00;
                               char33_0[50] <= 32'h00003F00;
                               char33_0[51] <= 32'h00007F80;
                               char33_0[52] <= 32'h000FFFFC;
                               char33_0[53] <= 32'h000FFFFC;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//4
                           4'd5: begin
                               char33_0[  0] <= 32'h00000000;
                               char33_0[  1] <= 32'h00000000;
                               char33_0[  2] <= 32'h00000000;
                               char33_0[  3] <= 32'h00000000;
                               char33_0[  4] <= 32'h00000000;
                               char33_0[  5] <= 32'h00000000;
                               char33_0[  6] <= 32'h00000000;
                               char33_0[  7] <= 32'h00000000;
                               char33_0[  8] <= 32'h00000000;
                               char33_0[  9] <= 32'h00000000;
                               char33_0[10] <= 32'h00000000;
                               char33_0[11] <= 32'h03FFFFF0;
                               char33_0[12] <= 32'h03FFFFF0;
                               char33_0[13] <= 32'h03FFFFF0;
                               char33_0[14] <= 32'h03FFFFE0;
                               char33_0[15] <= 32'h03800000;
                               char33_0[16] <= 32'h03800000;
                               char33_0[17] <= 32'h03800000;
                               char33_0[18] <= 32'h03800000;
                               char33_0[19] <= 32'h03800000;
                               char33_0[20] <= 32'h07800000;
                               char33_0[21] <= 32'h07800000;
                               char33_0[22] <= 32'h07800000;
                               char33_0[23] <= 32'h07800000;
                               char33_0[24] <= 32'h07800000;
                               char33_0[25] <= 32'h07800000;
                               char33_0[26] <= 32'h078FF800;
                               char33_0[27] <= 32'h073FFE00;
                               char33_0[28] <= 32'h077FFF80;
                               char33_0[29] <= 32'h07FC3F80;
                               char33_0[30] <= 32'h07E00FC0;
                               char33_0[31] <= 32'h07C007E0;
                               char33_0[32] <= 32'h078007E0;
                               char33_0[33] <= 32'h078003F0;
                               char33_0[34] <= 32'h000003F0;
                               char33_0[35] <= 32'h000001F0;
                               char33_0[36] <= 32'h000001F8;
                               char33_0[37] <= 32'h000001F8;
                               char33_0[38] <= 32'h000001F8;
                               char33_0[39] <= 32'h000001F8;
                               char33_0[40] <= 32'h000001F8;
                               char33_0[41] <= 32'h078001F8;
                               char33_0[42] <= 32'h0FC001F8;
                               char33_0[43] <= 32'h1FC001F0;
                               char33_0[44] <= 32'h1FC001F0;
                               char33_0[45] <= 32'h1FC003F0;
                               char33_0[46] <= 32'h1F8003F0;
                               char33_0[47] <= 32'h1F8003E0;
                               char33_0[48] <= 32'h0F8007E0;
                               char33_0[49] <= 32'h078007C0;
                               char33_0[50] <= 32'h07C01F80;
                               char33_0[51] <= 32'h03F83F00;
                               char33_0[52] <= 32'h00FFFE00;
                               char33_0[53] <= 32'h003FF800;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//5
                           4'd6: begin
                               char33_0[0] <= 32'h00000000;
                               char33_0[1] <= 32'h00000000;
                               char33_0[2] <= 32'h00000000;
                               char33_0[3] <= 32'h00000000;
                               char33_0[4] <= 32'h00000000;
                               char33_0[5] <= 32'h00000000;
                               char33_0[6] <= 32'h00000000;
                               char33_0[7] <= 32'h00000000;
                               char33_0[8] <= 32'h00000000;
                               char33_0[9] <= 32'h00000000;
                               char33_0[10] <= 32'h0007FE00;
                               char33_0[11] <= 32'h001FFF80;
                               char33_0[12] <= 32'h003F0FC0;
                               char33_0[13] <= 32'h007C07C0;
                               char33_0[14] <= 32'h00F807E0;
                               char33_0[15] <= 32'h01F007E0;
                               char33_0[16] <= 32'h03E007E0;
                               char33_0[17] <= 32'h03C007E0;
                               char33_0[18] <= 32'h07C003C0;
                               char33_0[19] <= 32'h07C00000;
                               char33_0[20] <= 32'h0FC00000;
                               char33_0[21] <= 32'h0F800000;
                               char33_0[22] <= 32'h0F800000;
                               char33_0[23] <= 32'h1F800000;
                               char33_0[24] <= 32'h1F800000;
                               char33_0[25] <= 32'h1F800000;
                               char33_0[26] <= 32'h1F87FE00;
                               char33_0[27] <= 32'h1F9FFF80;
                               char33_0[28] <= 32'h1FBFFFC0;
                               char33_0[29] <= 32'h3FFE1FC0;
                               char33_0[30] <= 32'h3FF807E0;
                               char33_0[31] <= 32'h3FE003F0;
                               char33_0[32] <= 32'h3FE003F0;
                               char33_0[33] <= 32'h3FC001F8;
                               char33_0[34] <= 32'h3F8001F8;
                               char33_0[35] <= 32'h3F8001F8;
                               char33_0[36] <= 32'h3F8000F8;
                               char33_0[37] <= 32'h3F8000F8;
                               char33_0[38] <= 32'h3F8000F8;
                               char33_0[39] <= 32'h1F8000F8;
                               char33_0[40] <= 32'h1F8000F8;
                               char33_0[41] <= 32'h1F8000F8;
                               char33_0[42] <= 32'h1F8000F8;
                               char33_0[43] <= 32'h1F8000F8;
                               char33_0[44] <= 32'h0FC001F8;
                               char33_0[45] <= 32'h0FC001F8;
                               char33_0[46] <= 32'h0FC001F0;
                               char33_0[47] <= 32'h07E001F0;
                               char33_0[48] <= 32'h03E003E0;
                               char33_0[49] <= 32'h03F003E0;
                               char33_0[50] <= 32'h01F807C0;
                               char33_0[51] <= 32'h00FE1F80;
                               char33_0[52] <= 32'h007FFE00;
                               char33_0[53] <= 32'h001FF800;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//6
                           4'd7: begin
                               char33_0[0] <= 32'h00000000;
                               char33_0[1] <= 32'h00000000;
                               char33_0[2] <= 32'h00000000;
                               char33_0[3] <= 32'h00000000;
                               char33_0[4] <= 32'h00000000;
                               char33_0[5] <= 32'h00000000;
                               char33_0[6] <= 32'h00000000;
                               char33_0[7] <= 32'h00000000;
                               char33_0[8] <= 32'h00000000;
                               char33_0[9] <= 32'h00000000;
                               char33_0[10] <= 32'h00000000;
                               char33_0[11] <= 32'h07FFFFF8;
                               char33_0[12] <= 32'h07FFFFF8;
                               char33_0[13] <= 32'h07FFFFF8;
                               char33_0[14] <= 32'h0FFFFFF0;
                               char33_0[15] <= 32'h0FC000E0;
                               char33_0[16] <= 32'h0F8001E0;
                               char33_0[17] <= 32'h0F0001C0;
                               char33_0[18] <= 32'h0E0003C0;
                               char33_0[19] <= 32'h0E000780;
                               char33_0[20] <= 32'h1E000780;
                               char33_0[21] <= 32'h1C000F00;
                               char33_0[22] <= 32'h00000F00;
                               char33_0[23] <= 32'h00001E00;
                               char33_0[24] <= 32'h00001E00;
                               char33_0[25] <= 32'h00003C00;
                               char33_0[26] <= 32'h00003C00;
                               char33_0[27] <= 32'h00007800;
                               char33_0[28] <= 32'h00007800;
                               char33_0[29] <= 32'h0000F800;
                               char33_0[30] <= 32'h0000F000;
                               char33_0[31] <= 32'h0001F000;
                               char33_0[32] <= 32'h0001E000;
                               char33_0[33] <= 32'h0003E000;
                               char33_0[34] <= 32'h0003E000;
                               char33_0[35] <= 32'h0003E000;
                               char33_0[36] <= 32'h0007C000;
                               char33_0[37] <= 32'h0007C000;
                               char33_0[38] <= 32'h0007C000;
                               char33_0[39] <= 32'h000FC000;
                               char33_0[40] <= 32'h000FC000;
                               char33_0[41] <= 32'h000FC000;
                               char33_0[42] <= 32'h000FC000;
                               char33_0[43] <= 32'h001FC000;
                               char33_0[44] <= 32'h001FC000;
                               char33_0[45] <= 32'h001FC000;
                               char33_0[46] <= 32'h001FC000;
                               char33_0[47] <= 32'h001FC000;
                               char33_0[48] <= 32'h001FC000;
                               char33_0[49] <= 32'h001FC000;
                               char33_0[50] <= 32'h001FC000;
                               char33_0[51] <= 32'h001FC000;
                               char33_0[52] <= 32'h001FC000;
                               char33_0[53] <= 32'h000F8000;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//7
                           4'd8: begin
                               char33_0[0] <= 32'h00000000;
                               char33_0[1] <= 32'h00000000;
                               char33_0[2] <= 32'h00000000;
                               char33_0[3] <= 32'h00000000;
                               char33_0[4] <= 32'h00000000;
                               char33_0[5] <= 32'h00000000;
                               char33_0[6] <= 32'h00000000;
                               char33_0[7] <= 32'h00000000;
                               char33_0[8] <= 32'h00000000;
                               char33_0[9] <= 32'h00000000;
                               char33_0[10] <= 32'h003FF800;
                               char33_0[11] <= 32'h00FFFE00;
                               char33_0[12] <= 32'h01F81F80;
                               char33_0[13] <= 32'h03E00FC0;
                               char33_0[14] <= 32'h07C003E0;
                               char33_0[15] <= 32'h0F8003E0;
                               char33_0[16] <= 32'h0F8001F0;
                               char33_0[17] <= 32'h1F0001F0;
                               char33_0[18] <= 32'h1F0001F0;
                               char33_0[19] <= 32'h1F0001F0;
                               char33_0[20] <= 32'h1F0001F0;
                               char33_0[21] <= 32'h1F0001F0;
                               char33_0[22] <= 32'h1F8001F0;
                               char33_0[23] <= 32'h1FC001F0;
                               char33_0[24] <= 32'h0FC001F0;
                               char33_0[25] <= 32'h0FF003E0;
                               char33_0[26] <= 32'h07F803C0;
                               char33_0[27] <= 32'h03FE0F80;
                               char33_0[28] <= 32'h01FF9F00;
                               char33_0[29] <= 32'h00FFFE00;
                               char33_0[30] <= 32'h003FF800;
                               char33_0[31] <= 32'h007FFC00;
                               char33_0[32] <= 32'h01F7FF00;
                               char33_0[33] <= 32'h03E1FF80;
                               char33_0[34] <= 32'h07C07FC0;
                               char33_0[35] <= 32'h0F801FE0;
                               char33_0[36] <= 32'h0F800FE0;
                               char33_0[37] <= 32'h1F0007F0;
                               char33_0[38] <= 32'h1F0003F0;
                               char33_0[39] <= 32'h3E0001F8;
                               char33_0[40] <= 32'h3E0001F8;
                               char33_0[41] <= 32'h3E0001F8;
                               char33_0[42] <= 32'h3E0000F8;
                               char33_0[43] <= 32'h3E0000F8;
                               char33_0[44] <= 32'h3E0000F8;
                               char33_0[45] <= 32'h3E0000F8;
                               char33_0[46] <= 32'h1F0001F0;
                               char33_0[47] <= 32'h1F0001F0;
                               char33_0[48] <= 32'h0F8003E0;
                               char33_0[49] <= 32'h0FC003E0;
                               char33_0[50] <= 32'h07E007C0;
                               char33_0[51] <= 32'h01F83F80;
                               char33_0[52] <= 32'h00FFFE00;
                               char33_0[53] <= 32'h003FF800;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//8
                           4'd9: begin
                               char33_0[0] <= 32'h00000000;
                               char33_0[1] <= 32'h00000000;
                               char33_0[2] <= 32'h00000000;
                               char33_0[3] <= 32'h00000000;
                               char33_0[4] <= 32'h00000000;
                               char33_0[5] <= 32'h00000000;
                               char33_0[6] <= 32'h00000000;
                               char33_0[7] <= 32'h00000000;
                               char33_0[8] <= 32'h00000000;
                               char33_0[9] <= 32'h00000000;
                               char33_0[10] <= 32'h003FF000;
                               char33_0[11] <= 32'h00FFFC00;
                               char33_0[12] <= 32'h01F83F00;
                               char33_0[13] <= 32'h03E01F80;
                               char33_0[14] <= 32'h07C00F80;
                               char33_0[15] <= 32'h0FC007C0;
                               char33_0[16] <= 32'h0F8003E0;
                               char33_0[17] <= 32'h1F8003E0;
                               char33_0[18] <= 32'h1F0003F0;
                               char33_0[19] <= 32'h1F0003F0;
                               char33_0[20] <= 32'h3F0001F0;
                               char33_0[21] <= 32'h3F0001F0;
                               char33_0[22] <= 32'h3F0001F8;
                               char33_0[23] <= 32'h3F0001F8;
                               char33_0[24] <= 32'h3F0001F8;
                               char33_0[25] <= 32'h3F0001F8;
                               char33_0[26] <= 32'h3F0001F8;
                               char33_0[27] <= 32'h3F0001F8;
                               char33_0[28] <= 32'h3F0003F8;
                               char33_0[29] <= 32'h1F8003F8;
                               char33_0[30] <= 32'h1F8007F8;
                               char33_0[31] <= 32'h1F800FF8;
                               char33_0[32] <= 32'h0FC01FF8;
                               char33_0[33] <= 32'h0FE03FF8;
                               char33_0[34] <= 32'h07F8FDF8;
                               char33_0[35] <= 32'h03FFF9F8;
                               char33_0[36] <= 32'h01FFF1F8;
                               char33_0[37] <= 32'h003F83F8;
                               char33_0[38] <= 32'h000003F0;
                               char33_0[39] <= 32'h000003F0;
                               char33_0[40] <= 32'h000003F0;
                               char33_0[41] <= 32'h000003F0;
                               char33_0[42] <= 32'h000007E0;
                               char33_0[43] <= 32'h000007E0;
                               char33_0[44] <= 32'h000007C0;
                               char33_0[45] <= 32'h03C007C0;
                               char33_0[46] <= 32'h07C00F80;
                               char33_0[47] <= 32'h0FE00F80;
                               char33_0[48] <= 32'h0FE01F00;
                               char33_0[49] <= 32'h0FE03E00;
                               char33_0[50] <= 32'h07E07E00;
                               char33_0[51] <= 32'h07F1F800;
                               char33_0[52] <= 32'h03FFF000;
                               char33_0[53] <= 32'h00FFC000;
                               char33_0[54] <= 32'h00000000;
                               char33_0[55] <= 32'h00000000;
                               char33_0[56] <= 32'h00000000;
                               char33_0[57] <= 32'h00000000;
                               char33_0[58] <= 32'h00000000;
                               char33_0[59] <= 32'h00000000;
                               char33_0[60] <= 32'h00000000;
                               char33_0[61] <= 32'h00000000;
                               char33_0[62] <= 32'h00000000;
                               char33_0[63] <= 32'h00000000;
                           end//9
                           default: begin
                               char33_0[0] <= char33_0[0];
                               char33_0[1] <= char33_0[1];
                               char33_0[2] <= char33_0[2];
                               char33_0[3] <= char33_0[3];
                               char33_0[4] <= char33_0[4];
                               char33_0[5] <= char33_0[5];
                               char33_0[6] <= char33_0[6];
                               char33_0[7] <= char33_0[7];
                               char33_0[8] <= char33_0[8];
                               char33_0[9] <= char33_0[9];
                               char33_0[10] <= char33_0[10];
                               char33_0[11] <= char33_0[11];
                               char33_0[12] <= char33_0[12];
                               char33_0[13] <= char33_0[13];
                               char33_0[14] <= char33_0[14];
                               char33_0[15] <= char33_0[15];
                               char33_0[16] <= char33_0[16];
                               char33_0[17] <= char33_0[17];
                               char33_0[18] <= char33_0[18];
                               char33_0[19] <= char33_0[19];
                               char33_0[20] <= char33_0[20];
                               char33_0[21] <= char33_0[21];
                               char33_0[22] <= char33_0[22];
                               char33_0[23] <= char33_0[23];
                               char33_0[24] <= char33_0[24];
                               char33_0[25] <= char33_0[25];
                               char33_0[26] <= char33_0[26];
                               char33_0[27] <= char33_0[27];
                               char33_0[28] <= char33_0[28];
                               char33_0[29] <= char33_0[29];
                               char33_0[30] <= char33_0[30];
                               char33_0[31] <= char33_0[31];
                               char33_0[32] <= char33_0[32];
                               char33_0[33] <= char33_0[33];
                               char33_0[34] <= char33_0[34];
                               char33_0[35] <= char33_0[35];
                               char33_0[36] <= char33_0[36];
                               char33_0[37] <= char33_0[37];
                               char33_0[38] <= char33_0[38];
                               char33_0[39] <= char33_0[39];
                               char33_0[40] <= char33_0[40];
                               char33_0[41] <= char33_0[41];
                               char33_0[42] <= char33_0[42];
                               char33_0[43] <= char33_0[43];
                               char33_0[44] <= char33_0[44];
                               char33_0[45] <= char33_0[45];
                               char33_0[46] <= char33_0[46];
                               char33_0[47] <= char33_0[47];
                               char33_0[48] <= char33_0[48];
                               char33_0[49] <= char33_0[49];
                               char33_0[50] <= char33_0[50];
                               char33_0[51] <= char33_0[51];
                               char33_0[52] <= char33_0[52];
                               char33_0[53] <= char33_0[53];
                               char33_0[54] <= char33_0[54];
                               char33_0[55] <= char33_0[55];
                               char33_0[56] <= char33_0[56];
                               char33_0[57] <= char33_0[57];
                               char33_0[58] <= char33_0[58];
                               char33_0[59] <= char33_0[59];
                               char33_0[60] <= char33_0[60];
                               char33_0[61] <= char33_0[61];
                               char33_0[62] <= char33_0[62];
                               char33_0[63] <= char33_0[63];
                           end
                       endcase
                   
                       case((a1 - w1*(a1/w1))/k1)
                               4'd0: begin
                                   char33_1[  0] <= 32'h00000000;
                                   char33_1[  1] <= 32'h00000000;
                                   char33_1[  2] <= 32'h00000000;
                                   char33_1[  3] <= 32'h00000000;
                                   char33_1[  4] <= 32'h00000000;
                                   char33_1[  5] <= 32'h00000000;
                                   char33_1[  6] <= 32'h00000000;
                                   char33_1[  7] <= 32'h00000000;
                                   char33_1[  8] <= 32'h00000000;
                                   char33_1[  9] <= 32'h00000000;
                                   char33_1[10] <= 32'h000FF000;
                                   char33_1[11] <= 32'h003FFC00;
                                   char33_1[12] <= 32'h007E7E00;
                                   char33_1[13] <= 32'h00F81F00;
                                   char33_1[14] <= 32'h01F00F80;
                                   char33_1[15] <= 32'h03F00FC0;
                                   char33_1[16] <= 32'h03E007C0;
                                   char33_1[17] <= 32'h07E007E0;
                                   char33_1[18] <= 32'h07C003E0;
                                   char33_1[19] <= 32'h0FC003F0;
                                   char33_1[20] <= 32'h0FC003F0;
                                   char33_1[21] <= 32'h0FC003F0;
                                   char33_1[22] <= 32'h1F8001F8;
                                   char33_1[23] <= 32'h1F8001F8;
                                   char33_1[24] <= 32'h1F8001F8;
                                   char33_1[25] <= 32'h1F8001F8;
                                   char33_1[26] <= 32'h1F8001F8;
                                   char33_1[27] <= 32'h3F8001F8;
                                   char33_1[28] <= 32'h3F8001F8;
                                   char33_1[29] <= 32'h3F8001F8;
                                   char33_1[30] <= 32'h3F8001F8;
                                   char33_1[31] <= 32'h3F8001F8;
                                   char33_1[32] <= 32'h3F8001F8;
                                   char33_1[33] <= 32'h3F8001F8;
                                   char33_1[34] <= 32'h3F8001F8;
                                   char33_1[35] <= 32'h3F8001F8;
                                   char33_1[36] <= 32'h3F8001F8;
                                   char33_1[37] <= 32'h1F8001F8;
                                   char33_1[38] <= 32'h1F8001F8;
                                   char33_1[39] <= 32'h1F8001F8;
                                   char33_1[40] <= 32'h1F8001F8;
                                   char33_1[41] <= 32'h1F8001F0;
                                   char33_1[42] <= 32'h0F8003F0;
                                   char33_1[43] <= 32'h0FC003F0;
                                   char33_1[44] <= 32'h0FC003F0;
                                   char33_1[45] <= 32'h07C003E0;
                                   char33_1[46] <= 32'h07E007E0;
                                   char33_1[47] <= 32'h03E007C0;
                                   char33_1[48] <= 32'h03F00FC0;
                                   char33_1[49] <= 32'h01F00F80;
                                   char33_1[50] <= 32'h00F81F00;
                                   char33_1[51] <= 32'h007E7E00;
                                   char33_1[52] <= 32'h003FFC00;
                                   char33_1[53] <= 32'h000FF000;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//0
                               4'd1: begin
                                   char33_1[  0] <= 32'h00000000;
                                   char33_1[  1] <= 32'h00000000;
                                   char33_1[  2] <= 32'h00000000;
                                   char33_1[  3] <= 32'h00000000;
                                   char33_1[  4] <= 32'h00000000;
                                   char33_1[  5] <= 32'h00000000;
                                   char33_1[  6] <= 32'h00000000;
                                   char33_1[  7] <= 32'h00000000;
                                   char33_1[  8] <= 32'h00000000;
                                   char33_1[  9] <= 32'h00000000;
                                   char33_1[10] <= 32'h0000E000;
                                   char33_1[11] <= 32'h0001E000;
                                   char33_1[12] <= 32'h0003E000;
                                   char33_1[13] <= 32'h001FE000;
                                   char33_1[14] <= 32'h03FFE000;
                                   char33_1[15] <= 32'h03FFE000;
                                   char33_1[16] <= 32'h0007E000;
                                   char33_1[17] <= 32'h0007E000;
                                   char33_1[18] <= 32'h0007E000;
                                   char33_1[19] <= 32'h0007E000;
                                   char33_1[20] <= 32'h0007E000;
                                   char33_1[21] <= 32'h0007E000;
                                   char33_1[22] <= 32'h0007E000;
                                   char33_1[23] <= 32'h0007E000;
                                   char33_1[24] <= 32'h0007E000;
                                   char33_1[25] <= 32'h0007E000;
                                   char33_1[26] <= 32'h0007E000;
                                   char33_1[27] <= 32'h0007E000;
                                   char33_1[28] <= 32'h0007E000;
                                   char33_1[29] <= 32'h0007E000;
                                   char33_1[30] <= 32'h0007E000;
                                   char33_1[31] <= 32'h0007E000;
                                   char33_1[32] <= 32'h0007E000;
                                   char33_1[33] <= 32'h0007E000;
                                   char33_1[34] <= 32'h0007E000;
                                   char33_1[35] <= 32'h0007E000;
                                   char33_1[36] <= 32'h0007E000;
                                   char33_1[37] <= 32'h0007E000;
                                   char33_1[38] <= 32'h0007E000;
                                   char33_1[39] <= 32'h0007E000;
                                   char33_1[40] <= 32'h0007E000;
                                   char33_1[41] <= 32'h0007E000;
                                   char33_1[42] <= 32'h0007E000;
                                   char33_1[43] <= 32'h0007E000;
                                   char33_1[44] <= 32'h0007E000;
                                   char33_1[45] <= 32'h0007E000;
                                   char33_1[46] <= 32'h0007E000;
                                   char33_1[47] <= 32'h0007E000;
                                   char33_1[48] <= 32'h0007E000;
                                   char33_1[49] <= 32'h0007E000;
                                   char33_1[50] <= 32'h0007E000;
                                   char33_1[51] <= 32'h000FF800;
                                   char33_1[52] <= 32'h03FFFFC0;
                                   char33_1[53] <= 32'h03FFFFC0;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//1
                               4'd2: begin
                                   char33_1[  0] <= 32'h00000000;
                                   char33_1[  1] <= 32'h00000000;
                                   char33_1[  2] <= 32'h00000000;
                                   char33_1[  3] <= 32'h00000000;
                                   char33_1[  4] <= 32'h00000000;
                                   char33_1[  5] <= 32'h00000000;
                                   char33_1[  6] <= 32'h00000000;
                                   char33_1[  7] <= 32'h00000000;
                                   char33_1[  8] <= 32'h00000000;
                                   char33_1[  9] <= 32'h00000000;
                                   char33_1[10] <= 32'h001FFC00;
                                   char33_1[11] <= 32'h007FFF00;
                                   char33_1[12] <= 32'h01F83F80;
                                   char33_1[13] <= 32'h03E00FC0;
                                   char33_1[14] <= 32'h07C007E0;
                                   char33_1[15] <= 32'h078007E0;
                                   char33_1[16] <= 32'h0F8003F0;
                                   char33_1[17] <= 32'h0F8003F0;
                                   char33_1[18] <= 32'h1F8003F0;
                                   char33_1[19] <= 32'h1F8003F0;
                                   char33_1[20] <= 32'h1FC003F0;
                                   char33_1[21] <= 32'h1FC003F0;
                                   char33_1[22] <= 32'h1FC003F0;
                                   char33_1[23] <= 32'h0FC003F0;
                                   char33_1[24] <= 32'h07C003F0;
                                   char33_1[25] <= 32'h000003E0;
                                   char33_1[26] <= 32'h000007E0;
                                   char33_1[27] <= 32'h000007E0;
                                   char33_1[28] <= 32'h00000FC0;
                                   char33_1[29] <= 32'h00000F80;
                                   char33_1[30] <= 32'h00001F80;
                                   char33_1[31] <= 32'h00003F00;
                                   char33_1[32] <= 32'h00003E00;
                                   char33_1[33] <= 32'h00007C00;
                                   char33_1[34] <= 32'h0000F800;
                                   char33_1[35] <= 32'h0001F000;
                                   char33_1[36] <= 32'h0003E000;
                                   char33_1[37] <= 32'h0007C000;
                                   char33_1[38] <= 32'h000F8000;
                                   char33_1[39] <= 32'h001F0000;
                                   char33_1[40] <= 32'h003E0000;
                                   char33_1[41] <= 32'h007C0000;
                                   char33_1[42] <= 32'h00F80000;
                                   char33_1[43] <= 32'h01F00038;
                                   char33_1[44] <= 32'h01E00038;
                                   char33_1[45] <= 32'h03C00070;
                                   char33_1[46] <= 32'h07800070;
                                   char33_1[47] <= 32'h0F8000F0;
                                   char33_1[48] <= 32'h0F0000F0;
                                   char33_1[49] <= 32'h1E0003F0;
                                   char33_1[50] <= 32'h3FFFFFF0;
                                   char33_1[51] <= 32'h3FFFFFF0;
                                   char33_1[52] <= 32'h3FFFFFE0;
                                   char33_1[53] <= 32'h3FFFFFE0;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//2
                               4'd3: begin
                                   char33_1[  0] <= 32'h00000000;
                                   char33_1[  1] <= 32'h00000000;
                                   char33_1[  2] <= 32'h00000000;
                                   char33_1[  3] <= 32'h00000000;
                                   char33_1[  4] <= 32'h00000000;
                                   char33_1[  5] <= 32'h00000000;
                                   char33_1[  6] <= 32'h00000000;
                                   char33_1[  7] <= 32'h00000000;
                                   char33_1[  8] <= 32'h00000000;
                                   char33_1[  9] <= 32'h00000000;
                                   char33_1[10] <= 32'h003FF000;
                                   char33_1[11] <= 32'h00FFFC00;
                                   char33_1[12] <= 32'h01F07E00;
                                   char33_1[13] <= 32'h03C03F00;
                                   char33_1[14] <= 32'h07801F80;
                                   char33_1[15] <= 32'h0F800FC0;
                                   char33_1[16] <= 32'h0F800FC0;
                                   char33_1[17] <= 32'h0F8007E0;
                                   char33_1[18] <= 32'h0FC007E0;
                                   char33_1[19] <= 32'h0FC007E0;
                                   char33_1[20] <= 32'h0FC007E0;
                                   char33_1[21] <= 32'h07C007E0;
                                   char33_1[22] <= 32'h000007E0;
                                   char33_1[23] <= 32'h000007E0;
                                   char33_1[24] <= 32'h000007C0;
                                   char33_1[25] <= 32'h00000FC0;
                                   char33_1[26] <= 32'h00000F80;
                                   char33_1[27] <= 32'h00001F00;
                                   char33_1[28] <= 32'h00007E00;
                                   char33_1[29] <= 32'h0003FC00;
                                   char33_1[30] <= 32'h001FF000;
                                   char33_1[31] <= 32'h001FFC00;
                                   char33_1[32] <= 32'h0000FF00;
                                   char33_1[33] <= 32'h00001F80;
                                   char33_1[34] <= 32'h00000FC0;
                                   char33_1[35] <= 32'h000007E0;
                                   char33_1[36] <= 32'h000003E0;
                                   char33_1[37] <= 32'h000003F0;
                                   char33_1[38] <= 32'h000003F0;
                                   char33_1[39] <= 32'h000001F0;
                                   char33_1[40] <= 32'h000001F8;
                                   char33_1[41] <= 32'h000001F8;
                                   char33_1[42] <= 32'h078001F8;
                                   char33_1[43] <= 32'h0FC001F8;
                                   char33_1[44] <= 32'h1FC001F8;
                                   char33_1[45] <= 32'h1FC003F0;
                                   char33_1[46] <= 32'h1FC003F0;
                                   char33_1[47] <= 32'h1FC003E0;
                                   char33_1[48] <= 32'h0F8007E0;
                                   char33_1[49] <= 32'h0F8007C0;
                                   char33_1[50] <= 32'h07C01F80;
                                   char33_1[51] <= 32'h03F07F00;
                                   char33_1[52] <= 32'h01FFFE00;
                                   char33_1[53] <= 32'h003FF000;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//3
                               4'd4: begin
                                   char33_1[  0] <= 32'h00000000;
                                   char33_1[  1] <= 32'h00000000;
                                   char33_1[  2] <= 32'h00000000;
                                   char33_1[  3] <= 32'h00000000;
                                   char33_1[  4] <= 32'h00000000;
                                   char33_1[  5] <= 32'h00000000;
                                   char33_1[  6] <= 32'h00000000;
                                   char33_1[  7] <= 32'h00000000;
                                   char33_1[  8] <= 32'h00000000;
                                   char33_1[  9] <= 32'h00000000;
                                   char33_1[10] <= 32'h00001F00;
                                   char33_1[11] <= 32'h00001F00;
                                   char33_1[12] <= 32'h00003F00;
                                   char33_1[13] <= 32'h00003F00;
                                   char33_1[14] <= 32'h00007F00;
                                   char33_1[15] <= 32'h0000FF00;
                                   char33_1[16] <= 32'h0000FF00;
                                   char33_1[17] <= 32'h0001FF00;
                                   char33_1[18] <= 32'h0003FF00;
                                   char33_1[19] <= 32'h0003BF00;
                                   char33_1[20] <= 32'h0007BF00;
                                   char33_1[21] <= 32'h00073F00;
                                   char33_1[22] <= 32'h000F3F00;
                                   char33_1[23] <= 32'h001E3F00;
                                   char33_1[24] <= 32'h001C3F00;
                                   char33_1[25] <= 32'h003C3F00;
                                   char33_1[26] <= 32'h00783F00;
                                   char33_1[27] <= 32'h00783F00;
                                   char33_1[28] <= 32'h00F03F00;
                                   char33_1[29] <= 32'h00E03F00;
                                   char33_1[30] <= 32'h01E03F00;
                                   char33_1[31] <= 32'h03C03F00;
                                   char33_1[32] <= 32'h03803F00;
                                   char33_1[33] <= 32'h07803F00;
                                   char33_1[34] <= 32'h0F003F00;
                                   char33_1[35] <= 32'h0F003F00;
                                   char33_1[36] <= 32'h1E003F00;
                                   char33_1[37] <= 32'h1C003F00;
                                   char33_1[38] <= 32'h3C003F00;
                                   char33_1[39] <= 32'h7FFFFFFE;
                                   char33_1[40] <= 32'h7FFFFFFE;
                                   char33_1[41] <= 32'h00003F00;
                                   char33_1[42] <= 32'h00003F00;
                                   char33_1[43] <= 32'h00003F00;
                                   char33_1[44] <= 32'h00003F00;
                                   char33_1[45] <= 32'h00003F00;
                                   char33_1[46] <= 32'h00003F00;
                                   char33_1[47] <= 32'h00003F00;
                                   char33_1[48] <= 32'h00003F00;
                                   char33_1[49] <= 32'h00003F00;
                                   char33_1[50] <= 32'h00003F00;
                                   char33_1[51] <= 32'h00007F80;
                                   char33_1[52] <= 32'h000FFFFC;
                                   char33_1[53] <= 32'h000FFFFC;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//4
                               4'd5: begin
                                   char33_1[  0] <= 32'h00000000;
                                   char33_1[  1] <= 32'h00000000;
                                   char33_1[  2] <= 32'h00000000;
                                   char33_1[  3] <= 32'h00000000;
                                   char33_1[  4] <= 32'h00000000;
                                   char33_1[  5] <= 32'h00000000;
                                   char33_1[  6] <= 32'h00000000;
                                   char33_1[  7] <= 32'h00000000;
                                   char33_1[  8] <= 32'h00000000;
                                   char33_1[  9] <= 32'h00000000;
                                   char33_1[10] <= 32'h00000000;
                                   char33_1[11] <= 32'h03FFFFF0;
                                   char33_1[12] <= 32'h03FFFFF0;
                                   char33_1[13] <= 32'h03FFFFF0;
                                   char33_1[14] <= 32'h03FFFFE0;
                                   char33_1[15] <= 32'h03800000;
                                   char33_1[16] <= 32'h03800000;
                                   char33_1[17] <= 32'h03800000;
                                   char33_1[18] <= 32'h03800000;
                                   char33_1[19] <= 32'h03800000;
                                   char33_1[20] <= 32'h07800000;
                                   char33_1[21] <= 32'h07800000;
                                   char33_1[22] <= 32'h07800000;
                                   char33_1[23] <= 32'h07800000;
                                   char33_1[24] <= 32'h07800000;
                                   char33_1[25] <= 32'h07800000;
                                   char33_1[26] <= 32'h078FF800;
                                   char33_1[27] <= 32'h073FFE00;
                                   char33_1[28] <= 32'h077FFF80;
                                   char33_1[29] <= 32'h07FC3F80;
                                   char33_1[30] <= 32'h07E00FC0;
                                   char33_1[31] <= 32'h07C007E0;
                                   char33_1[32] <= 32'h078007E0;
                                   char33_1[33] <= 32'h078003F0;
                                   char33_1[34] <= 32'h000003F0;
                                   char33_1[35] <= 32'h000001F0;
                                   char33_1[36] <= 32'h000001F8;
                                   char33_1[37] <= 32'h000001F8;
                                   char33_1[38] <= 32'h000001F8;
                                   char33_1[39] <= 32'h000001F8;
                                   char33_1[40] <= 32'h000001F8;
                                   char33_1[41] <= 32'h078001F8;
                                   char33_1[42] <= 32'h0FC001F8;
                                   char33_1[43] <= 32'h1FC001F0;
                                   char33_1[44] <= 32'h1FC001F0;
                                   char33_1[45] <= 32'h1FC003F0;
                                   char33_1[46] <= 32'h1F8003F0;
                                   char33_1[47] <= 32'h1F8003E0;
                                   char33_1[48] <= 32'h0F8007E0;
                                   char33_1[49] <= 32'h078007C0;
                                   char33_1[50] <= 32'h07C01F80;
                                   char33_1[51] <= 32'h03F83F00;
                                   char33_1[52] <= 32'h00FFFE00;
                                   char33_1[53] <= 32'h003FF800;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//5
                               4'd6: begin
                                   char33_1[0] <= 32'h00000000;
                                   char33_1[1] <= 32'h00000000;
                                   char33_1[2] <= 32'h00000000;
                                   char33_1[3] <= 32'h00000000;
                                   char33_1[4] <= 32'h00000000;
                                   char33_1[5] <= 32'h00000000;
                                   char33_1[6] <= 32'h00000000;
                                   char33_1[7] <= 32'h00000000;
                                   char33_1[8] <= 32'h00000000;
                                   char33_1[9] <= 32'h00000000;
                                   char33_1[10] <= 32'h0007FE00;
                                   char33_1[11] <= 32'h001FFF80;
                                   char33_1[12] <= 32'h003F0FC0;
                                   char33_1[13] <= 32'h007C07C0;
                                   char33_1[14] <= 32'h00F807E0;
                                   char33_1[15] <= 32'h01F007E0;
                                   char33_1[16] <= 32'h03E007E0;
                                   char33_1[17] <= 32'h03C007E0;
                                   char33_1[18] <= 32'h07C003C0;
                                   char33_1[19] <= 32'h07C00000;
                                   char33_1[20] <= 32'h0FC00000;
                                   char33_1[21] <= 32'h0F800000;
                                   char33_1[22] <= 32'h0F800000;
                                   char33_1[23] <= 32'h1F800000;
                                   char33_1[24] <= 32'h1F800000;
                                   char33_1[25] <= 32'h1F800000;
                                   char33_1[26] <= 32'h1F87FE00;
                                   char33_1[27] <= 32'h1F9FFF80;
                                   char33_1[28] <= 32'h1FBFFFC0;
                                   char33_1[29] <= 32'h3FFE1FC0;
                                   char33_1[30] <= 32'h3FF807E0;
                                   char33_1[31] <= 32'h3FE003F0;
                                   char33_1[32] <= 32'h3FE003F0;
                                   char33_1[33] <= 32'h3FC001F8;
                                   char33_1[34] <= 32'h3F8001F8;
                                   char33_1[35] <= 32'h3F8001F8;
                                   char33_1[36] <= 32'h3F8000F8;
                                   char33_1[37] <= 32'h3F8000F8;
                                   char33_1[38] <= 32'h3F8000F8;
                                   char33_1[39] <= 32'h1F8000F8;
                                   char33_1[40] <= 32'h1F8000F8;
                                   char33_1[41] <= 32'h1F8000F8;
                                   char33_1[42] <= 32'h1F8000F8;
                                   char33_1[43] <= 32'h1F8000F8;
                                   char33_1[44] <= 32'h0FC001F8;
                                   char33_1[45] <= 32'h0FC001F8;
                                   char33_1[46] <= 32'h0FC001F0;
                                   char33_1[47] <= 32'h07E001F0;
                                   char33_1[48] <= 32'h03E003E0;
                                   char33_1[49] <= 32'h03F003E0;
                                   char33_1[50] <= 32'h01F807C0;
                                   char33_1[51] <= 32'h00FE1F80;
                                   char33_1[52] <= 32'h007FFE00;
                                   char33_1[53] <= 32'h001FF800;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//6
                               4'd7: begin
                                   char33_1[0] <= 32'h00000000;
                                   char33_1[1] <= 32'h00000000;
                                   char33_1[2] <= 32'h00000000;
                                   char33_1[3] <= 32'h00000000;
                                   char33_1[4] <= 32'h00000000;
                                   char33_1[5] <= 32'h00000000;
                                   char33_1[6] <= 32'h00000000;
                                   char33_1[7] <= 32'h00000000;
                                   char33_1[8] <= 32'h00000000;
                                   char33_1[9] <= 32'h00000000;
                                   char33_1[10] <= 32'h00000000;
                                   char33_1[11] <= 32'h07FFFFF8;
                                   char33_1[12] <= 32'h07FFFFF8;
                                   char33_1[13] <= 32'h07FFFFF8;
                                   char33_1[14] <= 32'h0FFFFFF0;
                                   char33_1[15] <= 32'h0FC000E0;
                                   char33_1[16] <= 32'h0F8001E0;
                                   char33_1[17] <= 32'h0F0001C0;
                                   char33_1[18] <= 32'h0E0003C0;
                                   char33_1[19] <= 32'h0E000780;
                                   char33_1[20] <= 32'h1E000780;
                                   char33_1[21] <= 32'h1C000F00;
                                   char33_1[22] <= 32'h00000F00;
                                   char33_1[23] <= 32'h00001E00;
                                   char33_1[24] <= 32'h00001E00;
                                   char33_1[25] <= 32'h00003C00;
                                   char33_1[26] <= 32'h00003C00;
                                   char33_1[27] <= 32'h00007800;
                                   char33_1[28] <= 32'h00007800;
                                   char33_1[29] <= 32'h0000F800;
                                   char33_1[30] <= 32'h0000F000;
                                   char33_1[31] <= 32'h0001F000;
                                   char33_1[32] <= 32'h0001E000;
                                   char33_1[33] <= 32'h0003E000;
                                   char33_1[34] <= 32'h0003E000;
                                   char33_1[35] <= 32'h0003E000;
                                   char33_1[36] <= 32'h0007C000;
                                   char33_1[37] <= 32'h0007C000;
                                   char33_1[38] <= 32'h0007C000;
                                   char33_1[39] <= 32'h000FC000;
                                   char33_1[40] <= 32'h000FC000;
                                   char33_1[41] <= 32'h000FC000;
                                   char33_1[42] <= 32'h000FC000;
                                   char33_1[43] <= 32'h001FC000;
                                   char33_1[44] <= 32'h001FC000;
                                   char33_1[45] <= 32'h001FC000;
                                   char33_1[46] <= 32'h001FC000;
                                   char33_1[47] <= 32'h001FC000;
                                   char33_1[48] <= 32'h001FC000;
                                   char33_1[49] <= 32'h001FC000;
                                   char33_1[50] <= 32'h001FC000;
                                   char33_1[51] <= 32'h001FC000;
                                   char33_1[52] <= 32'h001FC000;
                                   char33_1[53] <= 32'h000F8000;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//7
                               4'd8: begin
                                   char33_1[0] <= 32'h00000000;
                                   char33_1[1] <= 32'h00000000;
                                   char33_1[2] <= 32'h00000000;
                                   char33_1[3] <= 32'h00000000;
                                   char33_1[4] <= 32'h00000000;
                                   char33_1[5] <= 32'h00000000;
                                   char33_1[6] <= 32'h00000000;
                                   char33_1[7] <= 32'h00000000;
                                   char33_1[8] <= 32'h00000000;
                                   char33_1[9] <= 32'h00000000;
                                   char33_1[10] <= 32'h003FF800;
                                   char33_1[11] <= 32'h00FFFE00;
                                   char33_1[12] <= 32'h01F81F80;
                                   char33_1[13] <= 32'h03E00FC0;
                                   char33_1[14] <= 32'h07C003E0;
                                   char33_1[15] <= 32'h0F8003E0;
                                   char33_1[16] <= 32'h0F8001F0;
                                   char33_1[17] <= 32'h1F0001F0;
                                   char33_1[18] <= 32'h1F0001F0;
                                   char33_1[19] <= 32'h1F0001F0;
                                   char33_1[20] <= 32'h1F0001F0;
                                   char33_1[21] <= 32'h1F0001F0;
                                   char33_1[22] <= 32'h1F8001F0;
                                   char33_1[23] <= 32'h1FC001F0;
                                   char33_1[24] <= 32'h0FC001F0;
                                   char33_1[25] <= 32'h0FF003E0;
                                   char33_1[26] <= 32'h07F803C0;
                                   char33_1[27] <= 32'h03FE0F80;
                                   char33_1[28] <= 32'h01FF9F00;
                                   char33_1[29] <= 32'h00FFFE00;
                                   char33_1[30] <= 32'h003FF800;
                                   char33_1[31] <= 32'h007FFC00;
                                   char33_1[32] <= 32'h01F7FF00;
                                   char33_1[33] <= 32'h03E1FF80;
                                   char33_1[34] <= 32'h07C07FC0;
                                   char33_1[35] <= 32'h0F801FE0;
                                   char33_1[36] <= 32'h0F800FE0;
                                   char33_1[37] <= 32'h1F0007F0;
                                   char33_1[38] <= 32'h1F0003F0;
                                   char33_1[39] <= 32'h3E0001F8;
                                   char33_1[40] <= 32'h3E0001F8;
                                   char33_1[41] <= 32'h3E0001F8;
                                   char33_1[42] <= 32'h3E0000F8;
                                   char33_1[43] <= 32'h3E0000F8;
                                   char33_1[44] <= 32'h3E0000F8;
                                   char33_1[45] <= 32'h3E0000F8;
                                   char33_1[46] <= 32'h1F0001F0;
                                   char33_1[47] <= 32'h1F0001F0;
                                   char33_1[48] <= 32'h0F8003E0;
                                   char33_1[49] <= 32'h0FC003E0;
                                   char33_1[50] <= 32'h07E007C0;
                                   char33_1[51] <= 32'h01F83F80;
                                   char33_1[52] <= 32'h00FFFE00;
                                   char33_1[53] <= 32'h003FF800;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//8
                               4'd9: begin
                                   char33_1[0] <= 32'h00000000;
                                   char33_1[1] <= 32'h00000000;
                                   char33_1[2] <= 32'h00000000;
                                   char33_1[3] <= 32'h00000000;
                                   char33_1[4] <= 32'h00000000;
                                   char33_1[5] <= 32'h00000000;
                                   char33_1[6] <= 32'h00000000;
                                   char33_1[7] <= 32'h00000000;
                                   char33_1[8] <= 32'h00000000;
                                   char33_1[9] <= 32'h00000000;
                                   char33_1[10] <= 32'h003FF000;
                                   char33_1[11] <= 32'h00FFFC00;
                                   char33_1[12] <= 32'h01F83F00;
                                   char33_1[13] <= 32'h03E01F80;
                                   char33_1[14] <= 32'h07C00F80;
                                   char33_1[15] <= 32'h0FC007C0;
                                   char33_1[16] <= 32'h0F8003E0;
                                   char33_1[17] <= 32'h1F8003E0;
                                   char33_1[18] <= 32'h1F0003F0;
                                   char33_1[19] <= 32'h1F0003F0;
                                   char33_1[20] <= 32'h3F0001F0;
                                   char33_1[21] <= 32'h3F0001F0;
                                   char33_1[22] <= 32'h3F0001F8;
                                   char33_1[23] <= 32'h3F0001F8;
                                   char33_1[24] <= 32'h3F0001F8;
                                   char33_1[25] <= 32'h3F0001F8;
                                   char33_1[26] <= 32'h3F0001F8;
                                   char33_1[27] <= 32'h3F0001F8;
                                   char33_1[28] <= 32'h3F0003F8;
                                   char33_1[29] <= 32'h1F8003F8;
                                   char33_1[30] <= 32'h1F8007F8;
                                   char33_1[31] <= 32'h1F800FF8;
                                   char33_1[32] <= 32'h0FC01FF8;
                                   char33_1[33] <= 32'h0FE03FF8;
                                   char33_1[34] <= 32'h07F8FDF8;
                                   char33_1[35] <= 32'h03FFF9F8;
                                   char33_1[36] <= 32'h01FFF1F8;
                                   char33_1[37] <= 32'h003F83F8;
                                   char33_1[38] <= 32'h000003F0;
                                   char33_1[39] <= 32'h000003F0;
                                   char33_1[40] <= 32'h000003F0;
                                   char33_1[41] <= 32'h000003F0;
                                   char33_1[42] <= 32'h000007E0;
                                   char33_1[43] <= 32'h000007E0;
                                   char33_1[44] <= 32'h000007C0;
                                   char33_1[45] <= 32'h03C007C0;
                                   char33_1[46] <= 32'h07C00F80;
                                   char33_1[47] <= 32'h0FE00F80;
                                   char33_1[48] <= 32'h0FE01F00;
                                   char33_1[49] <= 32'h0FE03E00;
                                   char33_1[50] <= 32'h07E07E00;
                                   char33_1[51] <= 32'h07F1F800;
                                   char33_1[52] <= 32'h03FFF000;
                                   char33_1[53] <= 32'h00FFC000;
                                   char33_1[54] <= 32'h00000000;
                                   char33_1[55] <= 32'h00000000;
                                   char33_1[56] <= 32'h00000000;
                                   char33_1[57] <= 32'h00000000;
                                   char33_1[58] <= 32'h00000000;
                                   char33_1[59] <= 32'h00000000;
                                   char33_1[60] <= 32'h00000000;
                                   char33_1[61] <= 32'h00000000;
                                   char33_1[62] <= 32'h00000000;
                                   char33_1[63] <= 32'h00000000;
                               end//9
                               default: begin
                                   char33_1[0] <= char33_1[0];
                                   char33_1[1] <= char33_1[1];
                                   char33_1[2] <= char33_1[2];
                                   char33_1[3] <= char33_1[3];
                                   char33_1[4] <= char33_1[4];
                                   char33_1[5] <= char33_1[5];
                                   char33_1[6] <= char33_1[6];
                                   char33_1[7] <= char33_1[7];
                                   char33_1[8] <= char33_1[8];
                                   char33_1[9] <= char33_1[9];
                                   char33_1[10] <= char33_1[10];
                                   char33_1[11] <= char33_1[11];
                                   char33_1[12] <= char33_1[12];
                                   char33_1[13] <= char33_1[13];
                                   char33_1[14] <= char33_1[14];
                                   char33_1[15] <= char33_1[15];
                                   char33_1[16] <= char33_1[16];
                                   char33_1[17] <= char33_1[17];
                                   char33_1[18] <= char33_1[18];
                                   char33_1[19] <= char33_1[19];
                                   char33_1[20] <= char33_1[20];
                                   char33_1[21] <= char33_1[21];
                                   char33_1[22] <= char33_1[22];
                                   char33_1[23] <= char33_1[23];
                                   char33_1[24] <= char33_1[24];
                                   char33_1[25] <= char33_1[25];
                                   char33_1[26] <= char33_1[26];
                                   char33_1[27] <= char33_1[27];
                                   char33_1[28] <= char33_1[28];
                                   char33_1[29] <= char33_1[29];
                                   char33_1[30] <= char33_1[30];
                                   char33_1[31] <= char33_1[31];
                                   char33_1[32] <= char33_1[32];
                                   char33_1[33] <= char33_1[33];
                                   char33_1[34] <= char33_1[34];
                                   char33_1[35] <= char33_1[35];
                                   char33_1[36] <= char33_1[36];
                                   char33_1[37] <= char33_1[37];
                                   char33_1[38] <= char33_1[38];
                                   char33_1[39] <= char33_1[39];
                                   char33_1[40] <= char33_1[40];
                                   char33_1[41] <= char33_1[41];
                                   char33_1[42] <= char33_1[42];
                                   char33_1[43] <= char33_1[43];
                                   char33_1[44] <= char33_1[44];
                                   char33_1[45] <= char33_1[45];
                                   char33_1[46] <= char33_1[46];
                                   char33_1[47] <= char33_1[47];
                                   char33_1[48] <= char33_1[48];
                                   char33_1[49] <= char33_1[49];
                                   char33_1[50] <= char33_1[50];
                                   char33_1[51] <= char33_1[51];
                                   char33_1[52] <= char33_1[52];
                                   char33_1[53] <= char33_1[53];
                                   char33_1[54] <= char33_1[54];
                                   char33_1[55] <= char33_1[55];
                                   char33_1[56] <= char33_1[56];
                                   char33_1[57] <= char33_1[57];
                                   char33_1[58] <= char33_1[58];
                                   char33_1[59] <= char33_1[59];
                                   char33_1[60] <= char33_1[60];
                                   char33_1[61] <= char33_1[61];
                                   char33_1[62] <= char33_1[62];
                                   char33_1[63] <= char33_1[63];
                               end
                           endcase
                   
                       case((a1 - k1*(a1/k1))/h1)
                                   4'd0: begin
                                       char33_2[  0] <= 32'h00000000;
                                       char33_2[  1] <= 32'h00000000;
                                       char33_2[  2] <= 32'h00000000;
                                       char33_2[  3] <= 32'h00000000;
                                       char33_2[  4] <= 32'h00000000;
                                       char33_2[  5] <= 32'h00000000;
                                       char33_2[  6] <= 32'h00000000;
                                       char33_2[  7] <= 32'h00000000;
                                       char33_2[  8] <= 32'h00000000;
                                       char33_2[  9] <= 32'h00000000;
                                       char33_2[10] <= 32'h000FF000;
                                       char33_2[11] <= 32'h003FFC00;
                                       char33_2[12] <= 32'h007E7E00;
                                       char33_2[13] <= 32'h00F81F00;
                                       char33_2[14] <= 32'h01F00F80;
                                       char33_2[15] <= 32'h03F00FC0;
                                       char33_2[16] <= 32'h03E007C0;
                                       char33_2[17] <= 32'h07E007E0;
                                       char33_2[18] <= 32'h07C003E0;
                                       char33_2[19] <= 32'h0FC003F0;
                                       char33_2[20] <= 32'h0FC003F0;
                                       char33_2[21] <= 32'h0FC003F0;
                                       char33_2[22] <= 32'h1F8001F8;
                                       char33_2[23] <= 32'h1F8001F8;
                                       char33_2[24] <= 32'h1F8001F8;
                                       char33_2[25] <= 32'h1F8001F8;
                                       char33_2[26] <= 32'h1F8001F8;
                                       char33_2[27] <= 32'h3F8001F8;
                                       char33_2[28] <= 32'h3F8001F8;
                                       char33_2[29] <= 32'h3F8001F8;
                                       char33_2[30] <= 32'h3F8001F8;
                                       char33_2[31] <= 32'h3F8001F8;
                                       char33_2[32] <= 32'h3F8001F8;
                                       char33_2[33] <= 32'h3F8001F8;
                                       char33_2[34] <= 32'h3F8001F8;
                                       char33_2[35] <= 32'h3F8001F8;
                                       char33_2[36] <= 32'h3F8001F8;
                                       char33_2[37] <= 32'h1F8001F8;
                                       char33_2[38] <= 32'h1F8001F8;
                                       char33_2[39] <= 32'h1F8001F8;
                                       char33_2[40] <= 32'h1F8001F8;
                                       char33_2[41] <= 32'h1F8001F0;
                                       char33_2[42] <= 32'h0F8003F0;
                                       char33_2[43] <= 32'h0FC003F0;
                                       char33_2[44] <= 32'h0FC003F0;
                                       char33_2[45] <= 32'h07C003E0;
                                       char33_2[46] <= 32'h07E007E0;
                                       char33_2[47] <= 32'h03E007C0;
                                       char33_2[48] <= 32'h03F00FC0;
                                       char33_2[49] <= 32'h01F00F80;
                                       char33_2[50] <= 32'h00F81F00;
                                       char33_2[51] <= 32'h007E7E00;
                                       char33_2[52] <= 32'h003FFC00;
                                       char33_2[53] <= 32'h000FF000;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//0
                                   4'd1: begin
                                       char33_2[  0] <= 32'h00000000;
                                       char33_2[  1] <= 32'h00000000;
                                       char33_2[  2] <= 32'h00000000;
                                       char33_2[  3] <= 32'h00000000;
                                       char33_2[  4] <= 32'h00000000;
                                       char33_2[  5] <= 32'h00000000;
                                       char33_2[  6] <= 32'h00000000;
                                       char33_2[  7] <= 32'h00000000;
                                       char33_2[  8] <= 32'h00000000;
                                       char33_2[  9] <= 32'h00000000;
                                       char33_2[10] <= 32'h0000E000;
                                       char33_2[11] <= 32'h0001E000;
                                       char33_2[12] <= 32'h0003E000;
                                       char33_2[13] <= 32'h001FE000;
                                       char33_2[14] <= 32'h03FFE000;
                                       char33_2[15] <= 32'h03FFE000;
                                       char33_2[16] <= 32'h0007E000;
                                       char33_2[17] <= 32'h0007E000;
                                       char33_2[18] <= 32'h0007E000;
                                       char33_2[19] <= 32'h0007E000;
                                       char33_2[20] <= 32'h0007E000;
                                       char33_2[21] <= 32'h0007E000;
                                       char33_2[22] <= 32'h0007E000;
                                       char33_2[23] <= 32'h0007E000;
                                       char33_2[24] <= 32'h0007E000;
                                       char33_2[25] <= 32'h0007E000;
                                       char33_2[26] <= 32'h0007E000;
                                       char33_2[27] <= 32'h0007E000;
                                       char33_2[28] <= 32'h0007E000;
                                       char33_2[29] <= 32'h0007E000;
                                       char33_2[30] <= 32'h0007E000;
                                       char33_2[31] <= 32'h0007E000;
                                       char33_2[32] <= 32'h0007E000;
                                       char33_2[33] <= 32'h0007E000;
                                       char33_2[34] <= 32'h0007E000;
                                       char33_2[35] <= 32'h0007E000;
                                       char33_2[36] <= 32'h0007E000;
                                       char33_2[37] <= 32'h0007E000;
                                       char33_2[38] <= 32'h0007E000;
                                       char33_2[39] <= 32'h0007E000;
                                       char33_2[40] <= 32'h0007E000;
                                       char33_2[41] <= 32'h0007E000;
                                       char33_2[42] <= 32'h0007E000;
                                       char33_2[43] <= 32'h0007E000;
                                       char33_2[44] <= 32'h0007E000;
                                       char33_2[45] <= 32'h0007E000;
                                       char33_2[46] <= 32'h0007E000;
                                       char33_2[47] <= 32'h0007E000;
                                       char33_2[48] <= 32'h0007E000;
                                       char33_2[49] <= 32'h0007E000;
                                       char33_2[50] <= 32'h0007E000;
                                       char33_2[51] <= 32'h000FF800;
                                       char33_2[52] <= 32'h03FFFFC0;
                                       char33_2[53] <= 32'h03FFFFC0;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//1
                                   4'd2: begin
                                       char33_2[  0] <= 32'h00000000;
                                       char33_2[  1] <= 32'h00000000;
                                       char33_2[  2] <= 32'h00000000;
                                       char33_2[  3] <= 32'h00000000;
                                       char33_2[  4] <= 32'h00000000;
                                       char33_2[  5] <= 32'h00000000;
                                       char33_2[  6] <= 32'h00000000;
                                       char33_2[  7] <= 32'h00000000;
                                       char33_2[  8] <= 32'h00000000;
                                       char33_2[  9] <= 32'h00000000;
                                       char33_2[10] <= 32'h001FFC00;
                                       char33_2[11] <= 32'h007FFF00;
                                       char33_2[12] <= 32'h01F83F80;
                                       char33_2[13] <= 32'h03E00FC0;
                                       char33_2[14] <= 32'h07C007E0;
                                       char33_2[15] <= 32'h078007E0;
                                       char33_2[16] <= 32'h0F8003F0;
                                       char33_2[17] <= 32'h0F8003F0;
                                       char33_2[18] <= 32'h1F8003F0;
                                       char33_2[19] <= 32'h1F8003F0;
                                       char33_2[20] <= 32'h1FC003F0;
                                       char33_2[21] <= 32'h1FC003F0;
                                       char33_2[22] <= 32'h1FC003F0;
                                       char33_2[23] <= 32'h0FC003F0;
                                       char33_2[24] <= 32'h07C003F0;
                                       char33_2[25] <= 32'h000003E0;
                                       char33_2[26] <= 32'h000007E0;
                                       char33_2[27] <= 32'h000007E0;
                                       char33_2[28] <= 32'h00000FC0;
                                       char33_2[29] <= 32'h00000F80;
                                       char33_2[30] <= 32'h00001F80;
                                       char33_2[31] <= 32'h00003F00;
                                       char33_2[32] <= 32'h00003E00;
                                       char33_2[33] <= 32'h00007C00;
                                       char33_2[34] <= 32'h0000F800;
                                       char33_2[35] <= 32'h0001F000;
                                       char33_2[36] <= 32'h0003E000;
                                       char33_2[37] <= 32'h0007C000;
                                       char33_2[38] <= 32'h000F8000;
                                       char33_2[39] <= 32'h001F0000;
                                       char33_2[40] <= 32'h003E0000;
                                       char33_2[41] <= 32'h007C0000;
                                       char33_2[42] <= 32'h00F80000;
                                       char33_2[43] <= 32'h01F00038;
                                       char33_2[44] <= 32'h01E00038;
                                       char33_2[45] <= 32'h03C00070;
                                       char33_2[46] <= 32'h07800070;
                                       char33_2[47] <= 32'h0F8000F0;
                                       char33_2[48] <= 32'h0F0000F0;
                                       char33_2[49] <= 32'h1E0003F0;
                                       char33_2[50] <= 32'h3FFFFFF0;
                                       char33_2[51] <= 32'h3FFFFFF0;
                                       char33_2[52] <= 32'h3FFFFFE0;
                                       char33_2[53] <= 32'h3FFFFFE0;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//2
                                   4'd3: begin
                                       char33_2[  0] <= 32'h00000000;
                                       char33_2[  1] <= 32'h00000000;
                                       char33_2[  2] <= 32'h00000000;
                                       char33_2[  3] <= 32'h00000000;
                                       char33_2[  4] <= 32'h00000000;
                                       char33_2[  5] <= 32'h00000000;
                                       char33_2[  6] <= 32'h00000000;
                                       char33_2[  7] <= 32'h00000000;
                                       char33_2[  8] <= 32'h00000000;
                                       char33_2[  9] <= 32'h00000000;
                                       char33_2[10] <= 32'h003FF000;
                                       char33_2[11] <= 32'h00FFFC00;
                                       char33_2[12] <= 32'h01F07E00;
                                       char33_2[13] <= 32'h03C03F00;
                                       char33_2[14] <= 32'h07801F80;
                                       char33_2[15] <= 32'h0F800FC0;
                                       char33_2[16] <= 32'h0F800FC0;
                                       char33_2[17] <= 32'h0F8007E0;
                                       char33_2[18] <= 32'h0FC007E0;
                                       char33_2[19] <= 32'h0FC007E0;
                                       char33_2[20] <= 32'h0FC007E0;
                                       char33_2[21] <= 32'h07C007E0;
                                       char33_2[22] <= 32'h000007E0;
                                       char33_2[23] <= 32'h000007E0;
                                       char33_2[24] <= 32'h000007C0;
                                       char33_2[25] <= 32'h00000FC0;
                                       char33_2[26] <= 32'h00000F80;
                                       char33_2[27] <= 32'h00001F00;
                                       char33_2[28] <= 32'h00007E00;
                                       char33_2[29] <= 32'h0003FC00;
                                       char33_2[30] <= 32'h001FF000;
                                       char33_2[31] <= 32'h001FFC00;
                                       char33_2[32] <= 32'h0000FF00;
                                       char33_2[33] <= 32'h00001F80;
                                       char33_2[34] <= 32'h00000FC0;
                                       char33_2[35] <= 32'h000007E0;
                                       char33_2[36] <= 32'h000003E0;
                                       char33_2[37] <= 32'h000003F0;
                                       char33_2[38] <= 32'h000003F0;
                                       char33_2[39] <= 32'h000001F0;
                                       char33_2[40] <= 32'h000001F8;
                                       char33_2[41] <= 32'h000001F8;
                                       char33_2[42] <= 32'h078001F8;
                                       char33_2[43] <= 32'h0FC001F8;
                                       char33_2[44] <= 32'h1FC001F8;
                                       char33_2[45] <= 32'h1FC003F0;
                                       char33_2[46] <= 32'h1FC003F0;
                                       char33_2[47] <= 32'h1FC003E0;
                                       char33_2[48] <= 32'h0F8007E0;
                                       char33_2[49] <= 32'h0F8007C0;
                                       char33_2[50] <= 32'h07C01F80;
                                       char33_2[51] <= 32'h03F07F00;
                                       char33_2[52] <= 32'h01FFFE00;
                                       char33_2[53] <= 32'h003FF000;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//3
                                   4'd4: begin
                                       char33_2[  0] <= 32'h00000000;
                                       char33_2[  1] <= 32'h00000000;
                                       char33_2[  2] <= 32'h00000000;
                                       char33_2[  3] <= 32'h00000000;
                                       char33_2[  4] <= 32'h00000000;
                                       char33_2[  5] <= 32'h00000000;
                                       char33_2[  6] <= 32'h00000000;
                                       char33_2[  7] <= 32'h00000000;
                                       char33_2[  8] <= 32'h00000000;
                                       char33_2[  9] <= 32'h00000000;
                                       char33_2[10] <= 32'h00001F00;
                                       char33_2[11] <= 32'h00001F00;
                                       char33_2[12] <= 32'h00003F00;
                                       char33_2[13] <= 32'h00003F00;
                                       char33_2[14] <= 32'h00007F00;
                                       char33_2[15] <= 32'h0000FF00;
                                       char33_2[16] <= 32'h0000FF00;
                                       char33_2[17] <= 32'h0001FF00;
                                       char33_2[18] <= 32'h0003FF00;
                                       char33_2[19] <= 32'h0003BF00;
                                       char33_2[20] <= 32'h0007BF00;
                                       char33_2[21] <= 32'h00073F00;
                                       char33_2[22] <= 32'h000F3F00;
                                       char33_2[23] <= 32'h001E3F00;
                                       char33_2[24] <= 32'h001C3F00;
                                       char33_2[25] <= 32'h003C3F00;
                                       char33_2[26] <= 32'h00783F00;
                                       char33_2[27] <= 32'h00783F00;
                                       char33_2[28] <= 32'h00F03F00;
                                       char33_2[29] <= 32'h00E03F00;
                                       char33_2[30] <= 32'h01E03F00;
                                       char33_2[31] <= 32'h03C03F00;
                                       char33_2[32] <= 32'h03803F00;
                                       char33_2[33] <= 32'h07803F00;
                                       char33_2[34] <= 32'h0F003F00;
                                       char33_2[35] <= 32'h0F003F00;
                                       char33_2[36] <= 32'h1E003F00;
                                       char33_2[37] <= 32'h1C003F00;
                                       char33_2[38] <= 32'h3C003F00;
                                       char33_2[39] <= 32'h7FFFFFFE;
                                       char33_2[40] <= 32'h7FFFFFFE;
                                       char33_2[41] <= 32'h00003F00;
                                       char33_2[42] <= 32'h00003F00;
                                       char33_2[43] <= 32'h00003F00;
                                       char33_2[44] <= 32'h00003F00;
                                       char33_2[45] <= 32'h00003F00;
                                       char33_2[46] <= 32'h00003F00;
                                       char33_2[47] <= 32'h00003F00;
                                       char33_2[48] <= 32'h00003F00;
                                       char33_2[49] <= 32'h00003F00;
                                       char33_2[50] <= 32'h00003F00;
                                       char33_2[51] <= 32'h00007F80;
                                       char33_2[52] <= 32'h000FFFFC;
                                       char33_2[53] <= 32'h000FFFFC;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//4
                                   4'd5: begin
                                       char33_2[  0] <= 32'h00000000;
                                       char33_2[  1] <= 32'h00000000;
                                       char33_2[  2] <= 32'h00000000;
                                       char33_2[  3] <= 32'h00000000;
                                       char33_2[  4] <= 32'h00000000;
                                       char33_2[  5] <= 32'h00000000;
                                       char33_2[  6] <= 32'h00000000;
                                       char33_2[  7] <= 32'h00000000;
                                       char33_2[  8] <= 32'h00000000;
                                       char33_2[  9] <= 32'h00000000;
                                       char33_2[10] <= 32'h00000000;
                                       char33_2[11] <= 32'h03FFFFF0;
                                       char33_2[12] <= 32'h03FFFFF0;
                                       char33_2[13] <= 32'h03FFFFF0;
                                       char33_2[14] <= 32'h03FFFFE0;
                                       char33_2[15] <= 32'h03800000;
                                       char33_2[16] <= 32'h03800000;
                                       char33_2[17] <= 32'h03800000;
                                       char33_2[18] <= 32'h03800000;
                                       char33_2[19] <= 32'h03800000;
                                       char33_2[20] <= 32'h07800000;
                                       char33_2[21] <= 32'h07800000;
                                       char33_2[22] <= 32'h07800000;
                                       char33_2[23] <= 32'h07800000;
                                       char33_2[24] <= 32'h07800000;
                                       char33_2[25] <= 32'h07800000;
                                       char33_2[26] <= 32'h078FF800;
                                       char33_2[27] <= 32'h073FFE00;
                                       char33_2[28] <= 32'h077FFF80;
                                       char33_2[29] <= 32'h07FC3F80;
                                       char33_2[30] <= 32'h07E00FC0;
                                       char33_2[31] <= 32'h07C007E0;
                                       char33_2[32] <= 32'h078007E0;
                                       char33_2[33] <= 32'h078003F0;
                                       char33_2[34] <= 32'h000003F0;
                                       char33_2[35] <= 32'h000001F0;
                                       char33_2[36] <= 32'h000001F8;
                                       char33_2[37] <= 32'h000001F8;
                                       char33_2[38] <= 32'h000001F8;
                                       char33_2[39] <= 32'h000001F8;
                                       char33_2[40] <= 32'h000001F8;
                                       char33_2[41] <= 32'h078001F8;
                                       char33_2[42] <= 32'h0FC001F8;
                                       char33_2[43] <= 32'h1FC001F0;
                                       char33_2[44] <= 32'h1FC001F0;
                                       char33_2[45] <= 32'h1FC003F0;
                                       char33_2[46] <= 32'h1F8003F0;
                                       char33_2[47] <= 32'h1F8003E0;
                                       char33_2[48] <= 32'h0F8007E0;
                                       char33_2[49] <= 32'h078007C0;
                                       char33_2[50] <= 32'h07C01F80;
                                       char33_2[51] <= 32'h03F83F00;
                                       char33_2[52] <= 32'h00FFFE00;
                                       char33_2[53] <= 32'h003FF800;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//5
                                   4'd6: begin
                                       char33_2[0] <= 32'h00000000;
                                       char33_2[1] <= 32'h00000000;
                                       char33_2[2] <= 32'h00000000;
                                       char33_2[3] <= 32'h00000000;
                                       char33_2[4] <= 32'h00000000;
                                       char33_2[5] <= 32'h00000000;
                                       char33_2[6] <= 32'h00000000;
                                       char33_2[7] <= 32'h00000000;
                                       char33_2[8] <= 32'h00000000;
                                       char33_2[9] <= 32'h00000000;
                                       char33_2[10] <= 32'h0007FE00;
                                       char33_2[11] <= 32'h001FFF80;
                                       char33_2[12] <= 32'h003F0FC0;
                                       char33_2[13] <= 32'h007C07C0;
                                       char33_2[14] <= 32'h00F807E0;
                                       char33_2[15] <= 32'h01F007E0;
                                       char33_2[16] <= 32'h03E007E0;
                                       char33_2[17] <= 32'h03C007E0;
                                       char33_2[18] <= 32'h07C003C0;
                                       char33_2[19] <= 32'h07C00000;
                                       char33_2[20] <= 32'h0FC00000;
                                       char33_2[21] <= 32'h0F800000;
                                       char33_2[22] <= 32'h0F800000;
                                       char33_2[23] <= 32'h1F800000;
                                       char33_2[24] <= 32'h1F800000;
                                       char33_2[25] <= 32'h1F800000;
                                       char33_2[26] <= 32'h1F87FE00;
                                       char33_2[27] <= 32'h1F9FFF80;
                                       char33_2[28] <= 32'h1FBFFFC0;
                                       char33_2[29] <= 32'h3FFE1FC0;
                                       char33_2[30] <= 32'h3FF807E0;
                                       char33_2[31] <= 32'h3FE003F0;
                                       char33_2[32] <= 32'h3FE003F0;
                                       char33_2[33] <= 32'h3FC001F8;
                                       char33_2[34] <= 32'h3F8001F8;
                                       char33_2[35] <= 32'h3F8001F8;
                                       char33_2[36] <= 32'h3F8000F8;
                                       char33_2[37] <= 32'h3F8000F8;
                                       char33_2[38] <= 32'h3F8000F8;
                                       char33_2[39] <= 32'h1F8000F8;
                                       char33_2[40] <= 32'h1F8000F8;
                                       char33_2[41] <= 32'h1F8000F8;
                                       char33_2[42] <= 32'h1F8000F8;
                                       char33_2[43] <= 32'h1F8000F8;
                                       char33_2[44] <= 32'h0FC001F8;
                                       char33_2[45] <= 32'h0FC001F8;
                                       char33_2[46] <= 32'h0FC001F0;
                                       char33_2[47] <= 32'h07E001F0;
                                       char33_2[48] <= 32'h03E003E0;
                                       char33_2[49] <= 32'h03F003E0;
                                       char33_2[50] <= 32'h01F807C0;
                                       char33_2[51] <= 32'h00FE1F80;
                                       char33_2[52] <= 32'h007FFE00;
                                       char33_2[53] <= 32'h001FF800;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//6
                                   4'd7: begin
                                       char33_2[0] <= 32'h00000000;
                                       char33_2[1] <= 32'h00000000;
                                       char33_2[2] <= 32'h00000000;
                                       char33_2[3] <= 32'h00000000;
                                       char33_2[4] <= 32'h00000000;
                                       char33_2[5] <= 32'h00000000;
                                       char33_2[6] <= 32'h00000000;
                                       char33_2[7] <= 32'h00000000;
                                       char33_2[8] <= 32'h00000000;
                                       char33_2[9] <= 32'h00000000;
                                       char33_2[10] <= 32'h00000000;
                                       char33_2[11] <= 32'h07FFFFF8;
                                       char33_2[12] <= 32'h07FFFFF8;
                                       char33_2[13] <= 32'h07FFFFF8;
                                       char33_2[14] <= 32'h0FFFFFF0;
                                       char33_2[15] <= 32'h0FC000E0;
                                       char33_2[16] <= 32'h0F8001E0;
                                       char33_2[17] <= 32'h0F0001C0;
                                       char33_2[18] <= 32'h0E0003C0;
                                       char33_2[19] <= 32'h0E000780;
                                       char33_2[20] <= 32'h1E000780;
                                       char33_2[21] <= 32'h1C000F00;
                                       char33_2[22] <= 32'h00000F00;
                                       char33_2[23] <= 32'h00001E00;
                                       char33_2[24] <= 32'h00001E00;
                                       char33_2[25] <= 32'h00003C00;
                                       char33_2[26] <= 32'h00003C00;
                                       char33_2[27] <= 32'h00007800;
                                       char33_2[28] <= 32'h00007800;
                                       char33_2[29] <= 32'h0000F800;
                                       char33_2[30] <= 32'h0000F000;
                                       char33_2[31] <= 32'h0001F000;
                                       char33_2[32] <= 32'h0001E000;
                                       char33_2[33] <= 32'h0003E000;
                                       char33_2[34] <= 32'h0003E000;
                                       char33_2[35] <= 32'h0003E000;
                                       char33_2[36] <= 32'h0007C000;
                                       char33_2[37] <= 32'h0007C000;
                                       char33_2[38] <= 32'h0007C000;
                                       char33_2[39] <= 32'h000FC000;
                                       char33_2[40] <= 32'h000FC000;
                                       char33_2[41] <= 32'h000FC000;
                                       char33_2[42] <= 32'h000FC000;
                                       char33_2[43] <= 32'h001FC000;
                                       char33_2[44] <= 32'h001FC000;
                                       char33_2[45] <= 32'h001FC000;
                                       char33_2[46] <= 32'h001FC000;
                                       char33_2[47] <= 32'h001FC000;
                                       char33_2[48] <= 32'h001FC000;
                                       char33_2[49] <= 32'h001FC000;
                                       char33_2[50] <= 32'h001FC000;
                                       char33_2[51] <= 32'h001FC000;
                                       char33_2[52] <= 32'h001FC000;
                                       char33_2[53] <= 32'h000F8000;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//7
                                   4'd8: begin
                                       char33_2[0] <= 32'h00000000;
                                       char33_2[1] <= 32'h00000000;
                                       char33_2[2] <= 32'h00000000;
                                       char33_2[3] <= 32'h00000000;
                                       char33_2[4] <= 32'h00000000;
                                       char33_2[5] <= 32'h00000000;
                                       char33_2[6] <= 32'h00000000;
                                       char33_2[7] <= 32'h00000000;
                                       char33_2[8] <= 32'h00000000;
                                       char33_2[9] <= 32'h00000000;
                                       char33_2[10] <= 32'h003FF800;
                                       char33_2[11] <= 32'h00FFFE00;
                                       char33_2[12] <= 32'h01F81F80;
                                       char33_2[13] <= 32'h03E00FC0;
                                       char33_2[14] <= 32'h07C003E0;
                                       char33_2[15] <= 32'h0F8003E0;
                                       char33_2[16] <= 32'h0F8001F0;
                                       char33_2[17] <= 32'h1F0001F0;
                                       char33_2[18] <= 32'h1F0001F0;
                                       char33_2[19] <= 32'h1F0001F0;
                                       char33_2[20] <= 32'h1F0001F0;
                                       char33_2[21] <= 32'h1F0001F0;
                                       char33_2[22] <= 32'h1F8001F0;
                                       char33_2[23] <= 32'h1FC001F0;
                                       char33_2[24] <= 32'h0FC001F0;
                                       char33_2[25] <= 32'h0FF003E0;
                                       char33_2[26] <= 32'h07F803C0;
                                       char33_2[27] <= 32'h03FE0F80;
                                       char33_2[28] <= 32'h01FF9F00;
                                       char33_2[29] <= 32'h00FFFE00;
                                       char33_2[30] <= 32'h003FF800;
                                       char33_2[31] <= 32'h007FFC00;
                                       char33_2[32] <= 32'h01F7FF00;
                                       char33_2[33] <= 32'h03E1FF80;
                                       char33_2[34] <= 32'h07C07FC0;
                                       char33_2[35] <= 32'h0F801FE0;
                                       char33_2[36] <= 32'h0F800FE0;
                                       char33_2[37] <= 32'h1F0007F0;
                                       char33_2[38] <= 32'h1F0003F0;
                                       char33_2[39] <= 32'h3E0001F8;
                                       char33_2[40] <= 32'h3E0001F8;
                                       char33_2[41] <= 32'h3E0001F8;
                                       char33_2[42] <= 32'h3E0000F8;
                                       char33_2[43] <= 32'h3E0000F8;
                                       char33_2[44] <= 32'h3E0000F8;
                                       char33_2[45] <= 32'h3E0000F8;
                                       char33_2[46] <= 32'h1F0001F0;
                                       char33_2[47] <= 32'h1F0001F0;
                                       char33_2[48] <= 32'h0F8003E0;
                                       char33_2[49] <= 32'h0FC003E0;
                                       char33_2[50] <= 32'h07E007C0;
                                       char33_2[51] <= 32'h01F83F80;
                                       char33_2[52] <= 32'h00FFFE00;
                                       char33_2[53] <= 32'h003FF800;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//8
                                   4'd9: begin
                                       char33_2[0] <= 32'h00000000;
                                       char33_2[1] <= 32'h00000000;
                                       char33_2[2] <= 32'h00000000;
                                       char33_2[3] <= 32'h00000000;
                                       char33_2[4] <= 32'h00000000;
                                       char33_2[5] <= 32'h00000000;
                                       char33_2[6] <= 32'h00000000;
                                       char33_2[7] <= 32'h00000000;
                                       char33_2[8] <= 32'h00000000;
                                       char33_2[9] <= 32'h00000000;
                                       char33_2[10] <= 32'h003FF000;
                                       char33_2[11] <= 32'h00FFFC00;
                                       char33_2[12] <= 32'h01F83F00;
                                       char33_2[13] <= 32'h03E01F80;
                                       char33_2[14] <= 32'h07C00F80;
                                       char33_2[15] <= 32'h0FC007C0;
                                       char33_2[16] <= 32'h0F8003E0;
                                       char33_2[17] <= 32'h1F8003E0;
                                       char33_2[18] <= 32'h1F0003F0;
                                       char33_2[19] <= 32'h1F0003F0;
                                       char33_2[20] <= 32'h3F0001F0;
                                       char33_2[21] <= 32'h3F0001F0;
                                       char33_2[22] <= 32'h3F0001F8;
                                       char33_2[23] <= 32'h3F0001F8;
                                       char33_2[24] <= 32'h3F0001F8;
                                       char33_2[25] <= 32'h3F0001F8;
                                       char33_2[26] <= 32'h3F0001F8;
                                       char33_2[27] <= 32'h3F0001F8;
                                       char33_2[28] <= 32'h3F0003F8;
                                       char33_2[29] <= 32'h1F8003F8;
                                       char33_2[30] <= 32'h1F8007F8;
                                       char33_2[31] <= 32'h1F800FF8;
                                       char33_2[32] <= 32'h0FC01FF8;
                                       char33_2[33] <= 32'h0FE03FF8;
                                       char33_2[34] <= 32'h07F8FDF8;
                                       char33_2[35] <= 32'h03FFF9F8;
                                       char33_2[36] <= 32'h01FFF1F8;
                                       char33_2[37] <= 32'h003F83F8;
                                       char33_2[38] <= 32'h000003F0;
                                       char33_2[39] <= 32'h000003F0;
                                       char33_2[40] <= 32'h000003F0;
                                       char33_2[41] <= 32'h000003F0;
                                       char33_2[42] <= 32'h000007E0;
                                       char33_2[43] <= 32'h000007E0;
                                       char33_2[44] <= 32'h000007C0;
                                       char33_2[45] <= 32'h03C007C0;
                                       char33_2[46] <= 32'h07C00F80;
                                       char33_2[47] <= 32'h0FE00F80;
                                       char33_2[48] <= 32'h0FE01F00;
                                       char33_2[49] <= 32'h0FE03E00;
                                       char33_2[50] <= 32'h07E07E00;
                                       char33_2[51] <= 32'h07F1F800;
                                       char33_2[52] <= 32'h03FFF000;
                                       char33_2[53] <= 32'h00FFC000;
                                       char33_2[54] <= 32'h00000000;
                                       char33_2[55] <= 32'h00000000;
                                       char33_2[56] <= 32'h00000000;
                                       char33_2[57] <= 32'h00000000;
                                       char33_2[58] <= 32'h00000000;
                                       char33_2[59] <= 32'h00000000;
                                       char33_2[60] <= 32'h00000000;
                                       char33_2[61] <= 32'h00000000;
                                       char33_2[62] <= 32'h00000000;
                                       char33_2[63] <= 32'h00000000;
                                   end//9
                                   default: begin
                                       char33_2[0] <= char33_2[0];
                                       char33_2[1] <= char33_2[1];
                                       char33_2[2] <= char33_2[2];
                                       char33_2[3] <= char33_2[3];
                                       char33_2[4] <= char33_2[4];
                                       char33_2[5] <= char33_2[5];
                                       char33_2[6] <= char33_2[6];
                                       char33_2[7] <= char33_2[7];
                                       char33_2[8] <= char33_2[8];
                                       char33_2[9] <= char33_2[9];
                                       char33_2[10] <= char33_2[10];
                                       char33_2[11] <= char33_2[11];
                                       char33_2[12] <= char33_2[12];
                                       char33_2[13] <= char33_2[13];
                                       char33_2[14] <= char33_2[14];
                                       char33_2[15] <= char33_2[15];
                                       char33_2[16] <= char33_2[16];
                                       char33_2[17] <= char33_2[17];
                                       char33_2[18] <= char33_2[18];
                                       char33_2[19] <= char33_2[19];
                                       char33_2[20] <= char33_2[20];
                                       char33_2[21] <= char33_2[21];
                                       char33_2[22] <= char33_2[22];
                                       char33_2[23] <= char33_2[23];
                                       char33_2[24] <= char33_2[24];
                                       char33_2[25] <= char33_2[25];
                                       char33_2[26] <= char33_2[26];
                                       char33_2[27] <= char33_2[27];
                                       char33_2[28] <= char33_2[28];
                                       char33_2[29] <= char33_2[29];
                                       char33_2[30] <= char33_2[30];
                                       char33_2[31] <= char33_2[31];
                                       char33_2[32] <= char33_2[32];
                                       char33_2[33] <= char33_2[33];
                                       char33_2[34] <= char33_2[34];
                                       char33_2[35] <= char33_2[35];
                                       char33_2[36] <= char33_2[36];
                                       char33_2[37] <= char33_2[37];
                                       char33_2[38] <= char33_2[38];
                                       char33_2[39] <= char33_2[39];
                                       char33_2[40] <= char33_2[40];
                                       char33_2[41] <= char33_2[41];
                                       char33_2[42] <= char33_2[42];
                                       char33_2[43] <= char33_2[43];
                                       char33_2[44] <= char33_2[44];
                                       char33_2[45] <= char33_2[45];
                                       char33_2[46] <= char33_2[46];
                                       char33_2[47] <= char33_2[47];
                                       char33_2[48] <= char33_2[48];
                                       char33_2[49] <= char33_2[49];
                                       char33_2[50] <= char33_2[50];
                                       char33_2[51] <= char33_2[51];
                                       char33_2[52] <= char33_2[52];
                                       char33_2[53] <= char33_2[53];
                                       char33_2[54] <= char33_2[54];
                                       char33_2[55] <= char33_2[55];
                                       char33_2[56] <= char33_2[56];
                                       char33_2[57] <= char33_2[57];
                                       char33_2[58] <= char33_2[58];
                                       char33_2[59] <= char33_2[59];
                                       char33_2[60] <= char33_2[60];
                                       char33_2[61] <= char33_2[61];
                                       char33_2[62] <= char33_2[62];
                                       char33_2[63] <= char33_2[63];
                                   end
                               endcase
                   
                        case((a1 - h1*(a1/h1))/t1)
                                       4'd0: begin
                                           char33_3[  0] <= 32'h00000000;
                                           char33_3[  1] <= 32'h00000000;
                                           char33_3[  2] <= 32'h00000000;
                                           char33_3[  3] <= 32'h00000000;
                                           char33_3[  4] <= 32'h00000000;
                                           char33_3[  5] <= 32'h00000000;
                                           char33_3[  6] <= 32'h00000000;
                                           char33_3[  7] <= 32'h00000000;
                                           char33_3[  8] <= 32'h00000000;
                                           char33_3[  9] <= 32'h00000000;
                                           char33_3[10] <= 32'h000FF000;
                                           char33_3[11] <= 32'h003FFC00;
                                           char33_3[12] <= 32'h007E7E00;
                                           char33_3[13] <= 32'h00F81F00;
                                           char33_3[14] <= 32'h01F00F80;
                                           char33_3[15] <= 32'h03F00FC0;
                                           char33_3[16] <= 32'h03E007C0;
                                           char33_3[17] <= 32'h07E007E0;
                                           char33_3[18] <= 32'h07C003E0;
                                           char33_3[19] <= 32'h0FC003F0;
                                           char33_3[20] <= 32'h0FC003F0;
                                           char33_3[21] <= 32'h0FC003F0;
                                           char33_3[22] <= 32'h1F8001F8;
                                           char33_3[23] <= 32'h1F8001F8;
                                           char33_3[24] <= 32'h1F8001F8;
                                           char33_3[25] <= 32'h1F8001F8;
                                           char33_3[26] <= 32'h1F8001F8;
                                           char33_3[27] <= 32'h3F8001F8;
                                           char33_3[28] <= 32'h3F8001F8;
                                           char33_3[29] <= 32'h3F8001F8;
                                           char33_3[30] <= 32'h3F8001F8;
                                           char33_3[31] <= 32'h3F8001F8;
                                           char33_3[32] <= 32'h3F8001F8;
                                           char33_3[33] <= 32'h3F8001F8;
                                           char33_3[34] <= 32'h3F8001F8;
                                           char33_3[35] <= 32'h3F8001F8;
                                           char33_3[36] <= 32'h3F8001F8;
                                           char33_3[37] <= 32'h1F8001F8;
                                           char33_3[38] <= 32'h1F8001F8;
                                           char33_3[39] <= 32'h1F8001F8;
                                           char33_3[40] <= 32'h1F8001F8;
                                           char33_3[41] <= 32'h1F8001F0;
                                           char33_3[42] <= 32'h0F8003F0;
                                           char33_3[43] <= 32'h0FC003F0;
                                           char33_3[44] <= 32'h0FC003F0;
                                           char33_3[45] <= 32'h07C003E0;
                                           char33_3[46] <= 32'h07E007E0;
                                           char33_3[47] <= 32'h03E007C0;
                                           char33_3[48] <= 32'h03F00FC0;
                                           char33_3[49] <= 32'h01F00F80;
                                           char33_3[50] <= 32'h00F81F00;
                                           char33_3[51] <= 32'h007E7E00;
                                           char33_3[52] <= 32'h003FFC00;
                                           char33_3[53] <= 32'h000FF000;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//0
                                       4'd1: begin
                                           char33_3[  0] <= 32'h00000000;
                                           char33_3[  1] <= 32'h00000000;
                                           char33_3[  2] <= 32'h00000000;
                                           char33_3[  3] <= 32'h00000000;
                                           char33_3[  4] <= 32'h00000000;
                                           char33_3[  5] <= 32'h00000000;
                                           char33_3[  6] <= 32'h00000000;
                                           char33_3[  7] <= 32'h00000000;
                                           char33_3[  8] <= 32'h00000000;
                                           char33_3[  9] <= 32'h00000000;
                                           char33_3[10] <= 32'h0000E000;
                                           char33_3[11] <= 32'h0001E000;
                                           char33_3[12] <= 32'h0003E000;
                                           char33_3[13] <= 32'h001FE000;
                                           char33_3[14] <= 32'h03FFE000;
                                           char33_3[15] <= 32'h03FFE000;
                                           char33_3[16] <= 32'h0007E000;
                                           char33_3[17] <= 32'h0007E000;
                                           char33_3[18] <= 32'h0007E000;
                                           char33_3[19] <= 32'h0007E000;
                                           char33_3[20] <= 32'h0007E000;
                                           char33_3[21] <= 32'h0007E000;
                                           char33_3[22] <= 32'h0007E000;
                                           char33_3[23] <= 32'h0007E000;
                                           char33_3[24] <= 32'h0007E000;
                                           char33_3[25] <= 32'h0007E000;
                                           char33_3[26] <= 32'h0007E000;
                                           char33_3[27] <= 32'h0007E000;
                                           char33_3[28] <= 32'h0007E000;
                                           char33_3[29] <= 32'h0007E000;
                                           char33_3[30] <= 32'h0007E000;
                                           char33_3[31] <= 32'h0007E000;
                                           char33_3[32] <= 32'h0007E000;
                                           char33_3[33] <= 32'h0007E000;
                                           char33_3[34] <= 32'h0007E000;
                                           char33_3[35] <= 32'h0007E000;
                                           char33_3[36] <= 32'h0007E000;
                                           char33_3[37] <= 32'h0007E000;
                                           char33_3[38] <= 32'h0007E000;
                                           char33_3[39] <= 32'h0007E000;
                                           char33_3[40] <= 32'h0007E000;
                                           char33_3[41] <= 32'h0007E000;
                                           char33_3[42] <= 32'h0007E000;
                                           char33_3[43] <= 32'h0007E000;
                                           char33_3[44] <= 32'h0007E000;
                                           char33_3[45] <= 32'h0007E000;
                                           char33_3[46] <= 32'h0007E000;
                                           char33_3[47] <= 32'h0007E000;
                                           char33_3[48] <= 32'h0007E000;
                                           char33_3[49] <= 32'h0007E000;
                                           char33_3[50] <= 32'h0007E000;
                                           char33_3[51] <= 32'h000FF800;
                                           char33_3[52] <= 32'h03FFFFC0;
                                           char33_3[53] <= 32'h03FFFFC0;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//1
                                       4'd2: begin
                                           char33_3[  0] <= 32'h00000000;
                                           char33_3[  1] <= 32'h00000000;
                                           char33_3[  2] <= 32'h00000000;
                                           char33_3[  3] <= 32'h00000000;
                                           char33_3[  4] <= 32'h00000000;
                                           char33_3[  5] <= 32'h00000000;
                                           char33_3[  6] <= 32'h00000000;
                                           char33_3[  7] <= 32'h00000000;
                                           char33_3[  8] <= 32'h00000000;
                                           char33_3[  9] <= 32'h00000000;
                                           char33_3[10] <= 32'h001FFC00;
                                           char33_3[11] <= 32'h007FFF00;
                                           char33_3[12] <= 32'h01F83F80;
                                           char33_3[13] <= 32'h03E00FC0;
                                           char33_3[14] <= 32'h07C007E0;
                                           char33_3[15] <= 32'h078007E0;
                                           char33_3[16] <= 32'h0F8003F0;
                                           char33_3[17] <= 32'h0F8003F0;
                                           char33_3[18] <= 32'h1F8003F0;
                                           char33_3[19] <= 32'h1F8003F0;
                                           char33_3[20] <= 32'h1FC003F0;
                                           char33_3[21] <= 32'h1FC003F0;
                                           char33_3[22] <= 32'h1FC003F0;
                                           char33_3[23] <= 32'h0FC003F0;
                                           char33_3[24] <= 32'h07C003F0;
                                           char33_3[25] <= 32'h000003E0;
                                           char33_3[26] <= 32'h000007E0;
                                           char33_3[27] <= 32'h000007E0;
                                           char33_3[28] <= 32'h00000FC0;
                                           char33_3[29] <= 32'h00000F80;
                                           char33_3[30] <= 32'h00001F80;
                                           char33_3[31] <= 32'h00003F00;
                                           char33_3[32] <= 32'h00003E00;
                                           char33_3[33] <= 32'h00007C00;
                                           char33_3[34] <= 32'h0000F800;
                                           char33_3[35] <= 32'h0001F000;
                                           char33_3[36] <= 32'h0003E000;
                                           char33_3[37] <= 32'h0007C000;
                                           char33_3[38] <= 32'h000F8000;
                                           char33_3[39] <= 32'h001F0000;
                                           char33_3[40] <= 32'h003E0000;
                                           char33_3[41] <= 32'h007C0000;
                                           char33_3[42] <= 32'h00F80000;
                                           char33_3[43] <= 32'h01F00038;
                                           char33_3[44] <= 32'h01E00038;
                                           char33_3[45] <= 32'h03C00070;
                                           char33_3[46] <= 32'h07800070;
                                           char33_3[47] <= 32'h0F8000F0;
                                           char33_3[48] <= 32'h0F0000F0;
                                           char33_3[49] <= 32'h1E0003F0;
                                           char33_3[50] <= 32'h3FFFFFF0;
                                           char33_3[51] <= 32'h3FFFFFF0;
                                           char33_3[52] <= 32'h3FFFFFE0;
                                           char33_3[53] <= 32'h3FFFFFE0;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//2
                                       4'd3: begin
                                           char33_3[  0] <= 32'h00000000;
                                           char33_3[  1] <= 32'h00000000;
                                           char33_3[  2] <= 32'h00000000;
                                           char33_3[  3] <= 32'h00000000;
                                           char33_3[  4] <= 32'h00000000;
                                           char33_3[  5] <= 32'h00000000;
                                           char33_3[  6] <= 32'h00000000;
                                           char33_3[  7] <= 32'h00000000;
                                           char33_3[  8] <= 32'h00000000;
                                           char33_3[  9] <= 32'h00000000;
                                           char33_3[10] <= 32'h003FF000;
                                           char33_3[11] <= 32'h00FFFC00;
                                           char33_3[12] <= 32'h01F07E00;
                                           char33_3[13] <= 32'h03C03F00;
                                           char33_3[14] <= 32'h07801F80;
                                           char33_3[15] <= 32'h0F800FC0;
                                           char33_3[16] <= 32'h0F800FC0;
                                           char33_3[17] <= 32'h0F8007E0;
                                           char33_3[18] <= 32'h0FC007E0;
                                           char33_3[19] <= 32'h0FC007E0;
                                           char33_3[20] <= 32'h0FC007E0;
                                           char33_3[21] <= 32'h07C007E0;
                                           char33_3[22] <= 32'h000007E0;
                                           char33_3[23] <= 32'h000007E0;
                                           char33_3[24] <= 32'h000007C0;
                                           char33_3[25] <= 32'h00000FC0;
                                           char33_3[26] <= 32'h00000F80;
                                           char33_3[27] <= 32'h00001F00;
                                           char33_3[28] <= 32'h00007E00;
                                           char33_3[29] <= 32'h0003FC00;
                                           char33_3[30] <= 32'h001FF000;
                                           char33_3[31] <= 32'h001FFC00;
                                           char33_3[32] <= 32'h0000FF00;
                                           char33_3[33] <= 32'h00001F80;
                                           char33_3[34] <= 32'h00000FC0;
                                           char33_3[35] <= 32'h000007E0;
                                           char33_3[36] <= 32'h000003E0;
                                           char33_3[37] <= 32'h000003F0;
                                           char33_3[38] <= 32'h000003F0;
                                           char33_3[39] <= 32'h000001F0;
                                           char33_3[40] <= 32'h000001F8;
                                           char33_3[41] <= 32'h000001F8;
                                           char33_3[42] <= 32'h078001F8;
                                           char33_3[43] <= 32'h0FC001F8;
                                           char33_3[44] <= 32'h1FC001F8;
                                           char33_3[45] <= 32'h1FC003F0;
                                           char33_3[46] <= 32'h1FC003F0;
                                           char33_3[47] <= 32'h1FC003E0;
                                           char33_3[48] <= 32'h0F8007E0;
                                           char33_3[49] <= 32'h0F8007C0;
                                           char33_3[50] <= 32'h07C01F80;
                                           char33_3[51] <= 32'h03F07F00;
                                           char33_3[52] <= 32'h01FFFE00;
                                           char33_3[53] <= 32'h003FF000;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//3
                                       4'd4: begin
                                           char33_3[  0] <= 32'h00000000;
                                           char33_3[  1] <= 32'h00000000;
                                           char33_3[  2] <= 32'h00000000;
                                           char33_3[  3] <= 32'h00000000;
                                           char33_3[  4] <= 32'h00000000;
                                           char33_3[  5] <= 32'h00000000;
                                           char33_3[  6] <= 32'h00000000;
                                           char33_3[  7] <= 32'h00000000;
                                           char33_3[  8] <= 32'h00000000;
                                           char33_3[  9] <= 32'h00000000;
                                           char33_3[10] <= 32'h00001F00;
                                           char33_3[11] <= 32'h00001F00;
                                           char33_3[12] <= 32'h00003F00;
                                           char33_3[13] <= 32'h00003F00;
                                           char33_3[14] <= 32'h00007F00;
                                           char33_3[15] <= 32'h0000FF00;
                                           char33_3[16] <= 32'h0000FF00;
                                           char33_3[17] <= 32'h0001FF00;
                                           char33_3[18] <= 32'h0003FF00;
                                           char33_3[19] <= 32'h0003BF00;
                                           char33_3[20] <= 32'h0007BF00;
                                           char33_3[21] <= 32'h00073F00;
                                           char33_3[22] <= 32'h000F3F00;
                                           char33_3[23] <= 32'h001E3F00;
                                           char33_3[24] <= 32'h001C3F00;
                                           char33_3[25] <= 32'h003C3F00;
                                           char33_3[26] <= 32'h00783F00;
                                           char33_3[27] <= 32'h00783F00;
                                           char33_3[28] <= 32'h00F03F00;
                                           char33_3[29] <= 32'h00E03F00;
                                           char33_3[30] <= 32'h01E03F00;
                                           char33_3[31] <= 32'h03C03F00;
                                           char33_3[32] <= 32'h03803F00;
                                           char33_3[33] <= 32'h07803F00;
                                           char33_3[34] <= 32'h0F003F00;
                                           char33_3[35] <= 32'h0F003F00;
                                           char33_3[36] <= 32'h1E003F00;
                                           char33_3[37] <= 32'h1C003F00;
                                           char33_3[38] <= 32'h3C003F00;
                                           char33_3[39] <= 32'h7FFFFFFE;
                                           char33_3[40] <= 32'h7FFFFFFE;
                                           char33_3[41] <= 32'h00003F00;
                                           char33_3[42] <= 32'h00003F00;
                                           char33_3[43] <= 32'h00003F00;
                                           char33_3[44] <= 32'h00003F00;
                                           char33_3[45] <= 32'h00003F00;
                                           char33_3[46] <= 32'h00003F00;
                                           char33_3[47] <= 32'h00003F00;
                                           char33_3[48] <= 32'h00003F00;
                                           char33_3[49] <= 32'h00003F00;
                                           char33_3[50] <= 32'h00003F00;
                                           char33_3[51] <= 32'h00007F80;
                                           char33_3[52] <= 32'h000FFFFC;
                                           char33_3[53] <= 32'h000FFFFC;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//4
                                       4'd5: begin
                                           char33_3[  0] <= 32'h00000000;
                                           char33_3[  1] <= 32'h00000000;
                                           char33_3[  2] <= 32'h00000000;
                                           char33_3[  3] <= 32'h00000000;
                                           char33_3[  4] <= 32'h00000000;
                                           char33_3[  5] <= 32'h00000000;
                                           char33_3[  6] <= 32'h00000000;
                                           char33_3[  7] <= 32'h00000000;
                                           char33_3[  8] <= 32'h00000000;
                                           char33_3[  9] <= 32'h00000000;
                                           char33_3[10] <= 32'h00000000;
                                           char33_3[11] <= 32'h03FFFFF0;
                                           char33_3[12] <= 32'h03FFFFF0;
                                           char33_3[13] <= 32'h03FFFFF0;
                                           char33_3[14] <= 32'h03FFFFE0;
                                           char33_3[15] <= 32'h03800000;
                                           char33_3[16] <= 32'h03800000;
                                           char33_3[17] <= 32'h03800000;
                                           char33_3[18] <= 32'h03800000;
                                           char33_3[19] <= 32'h03800000;
                                           char33_3[20] <= 32'h07800000;
                                           char33_3[21] <= 32'h07800000;
                                           char33_3[22] <= 32'h07800000;
                                           char33_3[23] <= 32'h07800000;
                                           char33_3[24] <= 32'h07800000;
                                           char33_3[25] <= 32'h07800000;
                                           char33_3[26] <= 32'h078FF800;
                                           char33_3[27] <= 32'h073FFE00;
                                           char33_3[28] <= 32'h077FFF80;
                                           char33_3[29] <= 32'h07FC3F80;
                                           char33_3[30] <= 32'h07E00FC0;
                                           char33_3[31] <= 32'h07C007E0;
                                           char33_3[32] <= 32'h078007E0;
                                           char33_3[33] <= 32'h078003F0;
                                           char33_3[34] <= 32'h000003F0;
                                           char33_3[35] <= 32'h000001F0;
                                           char33_3[36] <= 32'h000001F8;
                                           char33_3[37] <= 32'h000001F8;
                                           char33_3[38] <= 32'h000001F8;
                                           char33_3[39] <= 32'h000001F8;
                                           char33_3[40] <= 32'h000001F8;
                                           char33_3[41] <= 32'h078001F8;
                                           char33_3[42] <= 32'h0FC001F8;
                                           char33_3[43] <= 32'h1FC001F0;
                                           char33_3[44] <= 32'h1FC001F0;
                                           char33_3[45] <= 32'h1FC003F0;
                                           char33_3[46] <= 32'h1F8003F0;
                                           char33_3[47] <= 32'h1F8003E0;
                                           char33_3[48] <= 32'h0F8007E0;
                                           char33_3[49] <= 32'h078007C0;
                                           char33_3[50] <= 32'h07C01F80;
                                           char33_3[51] <= 32'h03F83F00;
                                           char33_3[52] <= 32'h00FFFE00;
                                           char33_3[53] <= 32'h003FF800;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//5
                                       4'd6: begin
                                           char33_3[0] <= 32'h00000000;
                                           char33_3[1] <= 32'h00000000;
                                           char33_3[2] <= 32'h00000000;
                                           char33_3[3] <= 32'h00000000;
                                           char33_3[4] <= 32'h00000000;
                                           char33_3[5] <= 32'h00000000;
                                           char33_3[6] <= 32'h00000000;
                                           char33_3[7] <= 32'h00000000;
                                           char33_3[8] <= 32'h00000000;
                                           char33_3[9] <= 32'h00000000;
                                           char33_3[10] <= 32'h0007FE00;
                                           char33_3[11] <= 32'h001FFF80;
                                           char33_3[12] <= 32'h003F0FC0;
                                           char33_3[13] <= 32'h007C07C0;
                                           char33_3[14] <= 32'h00F807E0;
                                           char33_3[15] <= 32'h01F007E0;
                                           char33_3[16] <= 32'h03E007E0;
                                           char33_3[17] <= 32'h03C007E0;
                                           char33_3[18] <= 32'h07C003C0;
                                           char33_3[19] <= 32'h07C00000;
                                           char33_3[20] <= 32'h0FC00000;
                                           char33_3[21] <= 32'h0F800000;
                                           char33_3[22] <= 32'h0F800000;
                                           char33_3[23] <= 32'h1F800000;
                                           char33_3[24] <= 32'h1F800000;
                                           char33_3[25] <= 32'h1F800000;
                                           char33_3[26] <= 32'h1F87FE00;
                                           char33_3[27] <= 32'h1F9FFF80;
                                           char33_3[28] <= 32'h1FBFFFC0;
                                           char33_3[29] <= 32'h3FFE1FC0;
                                           char33_3[30] <= 32'h3FF807E0;
                                           char33_3[31] <= 32'h3FE003F0;
                                           char33_3[32] <= 32'h3FE003F0;
                                           char33_3[33] <= 32'h3FC001F8;
                                           char33_3[34] <= 32'h3F8001F8;
                                           char33_3[35] <= 32'h3F8001F8;
                                           char33_3[36] <= 32'h3F8000F8;
                                           char33_3[37] <= 32'h3F8000F8;
                                           char33_3[38] <= 32'h3F8000F8;
                                           char33_3[39] <= 32'h1F8000F8;
                                           char33_3[40] <= 32'h1F8000F8;
                                           char33_3[41] <= 32'h1F8000F8;
                                           char33_3[42] <= 32'h1F8000F8;
                                           char33_3[43] <= 32'h1F8000F8;
                                           char33_3[44] <= 32'h0FC001F8;
                                           char33_3[45] <= 32'h0FC001F8;
                                           char33_3[46] <= 32'h0FC001F0;
                                           char33_3[47] <= 32'h07E001F0;
                                           char33_3[48] <= 32'h03E003E0;
                                           char33_3[49] <= 32'h03F003E0;
                                           char33_3[50] <= 32'h01F807C0;
                                           char33_3[51] <= 32'h00FE1F80;
                                           char33_3[52] <= 32'h007FFE00;
                                           char33_3[53] <= 32'h001FF800;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//6
                                       4'd7: begin
                                           char33_3[0] <= 32'h00000000;
                                           char33_3[1] <= 32'h00000000;
                                           char33_3[2] <= 32'h00000000;
                                           char33_3[3] <= 32'h00000000;
                                           char33_3[4] <= 32'h00000000;
                                           char33_3[5] <= 32'h00000000;
                                           char33_3[6] <= 32'h00000000;
                                           char33_3[7] <= 32'h00000000;
                                           char33_3[8] <= 32'h00000000;
                                           char33_3[9] <= 32'h00000000;
                                           char33_3[10] <= 32'h00000000;
                                           char33_3[11] <= 32'h07FFFFF8;
                                           char33_3[12] <= 32'h07FFFFF8;
                                           char33_3[13] <= 32'h07FFFFF8;
                                           char33_3[14] <= 32'h0FFFFFF0;
                                           char33_3[15] <= 32'h0FC000E0;
                                           char33_3[16] <= 32'h0F8001E0;
                                           char33_3[17] <= 32'h0F0001C0;
                                           char33_3[18] <= 32'h0E0003C0;
                                           char33_3[19] <= 32'h0E000780;
                                           char33_3[20] <= 32'h1E000780;
                                           char33_3[21] <= 32'h1C000F00;
                                           char33_3[22] <= 32'h00000F00;
                                           char33_3[23] <= 32'h00001E00;
                                           char33_3[24] <= 32'h00001E00;
                                           char33_3[25] <= 32'h00003C00;
                                           char33_3[26] <= 32'h00003C00;
                                           char33_3[27] <= 32'h00007800;
                                           char33_3[28] <= 32'h00007800;
                                           char33_3[29] <= 32'h0000F800;
                                           char33_3[30] <= 32'h0000F000;
                                           char33_3[31] <= 32'h0001F000;
                                           char33_3[32] <= 32'h0001E000;
                                           char33_3[33] <= 32'h0003E000;
                                           char33_3[34] <= 32'h0003E000;
                                           char33_3[35] <= 32'h0003E000;
                                           char33_3[36] <= 32'h0007C000;
                                           char33_3[37] <= 32'h0007C000;
                                           char33_3[38] <= 32'h0007C000;
                                           char33_3[39] <= 32'h000FC000;
                                           char33_3[40] <= 32'h000FC000;
                                           char33_3[41] <= 32'h000FC000;
                                           char33_3[42] <= 32'h000FC000;
                                           char33_3[43] <= 32'h001FC000;
                                           char33_3[44] <= 32'h001FC000;
                                           char33_3[45] <= 32'h001FC000;
                                           char33_3[46] <= 32'h001FC000;
                                           char33_3[47] <= 32'h001FC000;
                                           char33_3[48] <= 32'h001FC000;
                                           char33_3[49] <= 32'h001FC000;
                                           char33_3[50] <= 32'h001FC000;
                                           char33_3[51] <= 32'h001FC000;
                                           char33_3[52] <= 32'h001FC000;
                                           char33_3[53] <= 32'h000F8000;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//7
                                       4'd8: begin
                                           char33_3[0] <= 32'h00000000;
                                           char33_3[1] <= 32'h00000000;
                                           char33_3[2] <= 32'h00000000;
                                           char33_3[3] <= 32'h00000000;
                                           char33_3[4] <= 32'h00000000;
                                           char33_3[5] <= 32'h00000000;
                                           char33_3[6] <= 32'h00000000;
                                           char33_3[7] <= 32'h00000000;
                                           char33_3[8] <= 32'h00000000;
                                           char33_3[9] <= 32'h00000000;
                                           char33_3[10] <= 32'h003FF800;
                                           char33_3[11] <= 32'h00FFFE00;
                                           char33_3[12] <= 32'h01F81F80;
                                           char33_3[13] <= 32'h03E00FC0;
                                           char33_3[14] <= 32'h07C003E0;
                                           char33_3[15] <= 32'h0F8003E0;
                                           char33_3[16] <= 32'h0F8001F0;
                                           char33_3[17] <= 32'h1F0001F0;
                                           char33_3[18] <= 32'h1F0001F0;
                                           char33_3[19] <= 32'h1F0001F0;
                                           char33_3[20] <= 32'h1F0001F0;
                                           char33_3[21] <= 32'h1F0001F0;
                                           char33_3[22] <= 32'h1F8001F0;
                                           char33_3[23] <= 32'h1FC001F0;
                                           char33_3[24] <= 32'h0FC001F0;
                                           char33_3[25] <= 32'h0FF003E0;
                                           char33_3[26] <= 32'h07F803C0;
                                           char33_3[27] <= 32'h03FE0F80;
                                           char33_3[28] <= 32'h01FF9F00;
                                           char33_3[29] <= 32'h00FFFE00;
                                           char33_3[30] <= 32'h003FF800;
                                           char33_3[31] <= 32'h007FFC00;
                                           char33_3[32] <= 32'h01F7FF00;
                                           char33_3[33] <= 32'h03E1FF80;
                                           char33_3[34] <= 32'h07C07FC0;
                                           char33_3[35] <= 32'h0F801FE0;
                                           char33_3[36] <= 32'h0F800FE0;
                                           char33_3[37] <= 32'h1F0007F0;
                                           char33_3[38] <= 32'h1F0003F0;
                                           char33_3[39] <= 32'h3E0001F8;
                                           char33_3[40] <= 32'h3E0001F8;
                                           char33_3[41] <= 32'h3E0001F8;
                                           char33_3[42] <= 32'h3E0000F8;
                                           char33_3[43] <= 32'h3E0000F8;
                                           char33_3[44] <= 32'h3E0000F8;
                                           char33_3[45] <= 32'h3E0000F8;
                                           char33_3[46] <= 32'h1F0001F0;
                                           char33_3[47] <= 32'h1F0001F0;
                                           char33_3[48] <= 32'h0F8003E0;
                                           char33_3[49] <= 32'h0FC003E0;
                                           char33_3[50] <= 32'h07E007C0;
                                           char33_3[51] <= 32'h01F83F80;
                                           char33_3[52] <= 32'h00FFFE00;
                                           char33_3[53] <= 32'h003FF800;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//8
                                       4'd9: begin
                                           char33_3[0] <= 32'h00000000;
                                           char33_3[1] <= 32'h00000000;
                                           char33_3[2] <= 32'h00000000;
                                           char33_3[3] <= 32'h00000000;
                                           char33_3[4] <= 32'h00000000;
                                           char33_3[5] <= 32'h00000000;
                                           char33_3[6] <= 32'h00000000;
                                           char33_3[7] <= 32'h00000000;
                                           char33_3[8] <= 32'h00000000;
                                           char33_3[9] <= 32'h00000000;
                                           char33_3[10] <= 32'h003FF000;
                                           char33_3[11] <= 32'h00FFFC00;
                                           char33_3[12] <= 32'h01F83F00;
                                           char33_3[13] <= 32'h03E01F80;
                                           char33_3[14] <= 32'h07C00F80;
                                           char33_3[15] <= 32'h0FC007C0;
                                           char33_3[16] <= 32'h0F8003E0;
                                           char33_3[17] <= 32'h1F8003E0;
                                           char33_3[18] <= 32'h1F0003F0;
                                           char33_3[19] <= 32'h1F0003F0;
                                           char33_3[20] <= 32'h3F0001F0;
                                           char33_3[21] <= 32'h3F0001F0;
                                           char33_3[22] <= 32'h3F0001F8;
                                           char33_3[23] <= 32'h3F0001F8;
                                           char33_3[24] <= 32'h3F0001F8;
                                           char33_3[25] <= 32'h3F0001F8;
                                           char33_3[26] <= 32'h3F0001F8;
                                           char33_3[27] <= 32'h3F0001F8;
                                           char33_3[28] <= 32'h3F0003F8;
                                           char33_3[29] <= 32'h1F8003F8;
                                           char33_3[30] <= 32'h1F8007F8;
                                           char33_3[31] <= 32'h1F800FF8;
                                           char33_3[32] <= 32'h0FC01FF8;
                                           char33_3[33] <= 32'h0FE03FF8;
                                           char33_3[34] <= 32'h07F8FDF8;
                                           char33_3[35] <= 32'h03FFF9F8;
                                           char33_3[36] <= 32'h01FFF1F8;
                                           char33_3[37] <= 32'h003F83F8;
                                           char33_3[38] <= 32'h000003F0;
                                           char33_3[39] <= 32'h000003F0;
                                           char33_3[40] <= 32'h000003F0;
                                           char33_3[41] <= 32'h000003F0;
                                           char33_3[42] <= 32'h000007E0;
                                           char33_3[43] <= 32'h000007E0;
                                           char33_3[44] <= 32'h000007C0;
                                           char33_3[45] <= 32'h03C007C0;
                                           char33_3[46] <= 32'h07C00F80;
                                           char33_3[47] <= 32'h0FE00F80;
                                           char33_3[48] <= 32'h0FE01F00;
                                           char33_3[49] <= 32'h0FE03E00;
                                           char33_3[50] <= 32'h07E07E00;
                                           char33_3[51] <= 32'h07F1F800;
                                           char33_3[52] <= 32'h03FFF000;
                                           char33_3[53] <= 32'h00FFC000;
                                           char33_3[54] <= 32'h00000000;
                                           char33_3[55] <= 32'h00000000;
                                           char33_3[56] <= 32'h00000000;
                                           char33_3[57] <= 32'h00000000;
                                           char33_3[58] <= 32'h00000000;
                                           char33_3[59] <= 32'h00000000;
                                           char33_3[60] <= 32'h00000000;
                                           char33_3[61] <= 32'h00000000;
                                           char33_3[62] <= 32'h00000000;
                                           char33_3[63] <= 32'h00000000;
                                       end//9
                                       default: begin
                                           char33_3[0] <= char33_3[0];
                                           char33_3[1] <= char33_3[1];
                                           char33_3[2] <= char33_3[2];
                                           char33_3[3] <= char33_3[3];
                                           char33_3[4] <= char33_3[4];
                                           char33_3[5] <= char33_3[5];
                                           char33_3[6] <= char33_3[6];
                                           char33_3[7] <= char33_3[7];
                                           char33_3[8] <= char33_3[8];
                                           char33_3[9] <= char33_3[9];
                                           char33_3[10] <= char33_3[10];
                                           char33_3[11] <= char33_3[11];
                                           char33_3[12] <= char33_3[12];
                                           char33_3[13] <= char33_3[13];
                                           char33_3[14] <= char33_3[14];
                                           char33_3[15] <= char33_3[15];
                                           char33_3[16] <= char33_3[16];
                                           char33_3[17] <= char33_3[17];
                                           char33_3[18] <= char33_3[18];
                                           char33_3[19] <= char33_3[19];
                                           char33_3[20] <= char33_3[20];
                                           char33_3[21] <= char33_3[21];
                                           char33_3[22] <= char33_3[22];
                                           char33_3[23] <= char33_3[23];
                                           char33_3[24] <= char33_3[24];
                                           char33_3[25] <= char33_3[25];
                                           char33_3[26] <= char33_3[26];
                                           char33_3[27] <= char33_3[27];
                                           char33_3[28] <= char33_3[28];
                                           char33_3[29] <= char33_3[29];
                                           char33_3[30] <= char33_3[30];
                                           char33_3[31] <= char33_3[31];
                                           char33_3[32] <= char33_3[32];
                                           char33_3[33] <= char33_3[33];
                                           char33_3[34] <= char33_3[34];
                                           char33_3[35] <= char33_3[35];
                                           char33_3[36] <= char33_3[36];
                                           char33_3[37] <= char33_3[37];
                                           char33_3[38] <= char33_3[38];
                                           char33_3[39] <= char33_3[39];
                                           char33_3[40] <= char33_3[40];
                                           char33_3[41] <= char33_3[41];
                                           char33_3[42] <= char33_3[42];
                                           char33_3[43] <= char33_3[43];
                                           char33_3[44] <= char33_3[44];
                                           char33_3[45] <= char33_3[45];
                                           char33_3[46] <= char33_3[46];
                                           char33_3[47] <= char33_3[47];
                                           char33_3[48] <= char33_3[48];
                                           char33_3[49] <= char33_3[49];
                                           char33_3[50] <= char33_3[50];
                                           char33_3[51] <= char33_3[51];
                                           char33_3[52] <= char33_3[52];
                                           char33_3[53] <= char33_3[53];
                                           char33_3[54] <= char33_3[54];
                                           char33_3[55] <= char33_3[55];
                                           char33_3[56] <= char33_3[56];
                                           char33_3[57] <= char33_3[57];
                                           char33_3[58] <= char33_3[58];
                                           char33_3[59] <= char33_3[59];
                                           char33_3[60] <= char33_3[60];
                                           char33_3[61] <= char33_3[61];
                                           char33_3[62] <= char33_3[62];
                                           char33_3[63] <= char33_3[63];
                                       end
                                   endcase
                  
                       case((a1 - t1*(a1/t1))/o1)
                                  4'd0: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h000FF000000000000000000000000000;
                                        char33_4[11] <= 128'h003FFC00000000000000000000000000;
                                        char33_4[12] <= 128'h007E7E00800000000000000000000000;
                                        char33_4[13] <= 128'h00F81F00000000000000000000000000;
                                        char33_4[14] <= 128'h01F00F80000000000000000000000000;
                                        char33_4[15] <= 128'h03F00FC0000000000000000000000000;
                                        char33_4[16] <= 128'h03E007C0000000000000000000000000;
                                        char33_4[17] <= 128'h07E007E0000000000000000000000000;
                                        char33_4[18] <= 128'h07C003E0000000000000000000000000;
                                        char33_4[19] <= 128'h0FC003F0000000000000000000000000;
                                        char33_4[20] <= 128'h0FC003F0000000000000000000000000;
                                        char33_4[21] <= 128'h0FC003F0000000000000000000000000;
                                        char33_4[22] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[23] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[24] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[25] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[26] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[27] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[28] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[29] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[30] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[31] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[32] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[33] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[34] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[35] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[36] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[37] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[38] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[39] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[40] <= 128'h1F8001F8000000000000000000000000;
                                        char33_4[41] <= 128'h1F8001F0000000000000000000000000;
                                        char33_4[42] <= 128'h0F8003F0000000000000000000000000;
                                        char33_4[43] <= 128'h0FC003F0000000000000000000000000;
                                        char33_4[44] <= 128'h0FC003F0000000000000000000000000;
                                        char33_4[45] <= 128'h07C003E0000000000000000000000000;
                                        char33_4[46] <= 128'h07E007E0000000000000000000000000;
                                        char33_4[47] <= 128'h03E007C0000000000000000000000000;
                                        char33_4[48] <= 128'h03F00FC0000000000000000000000000;
                                        char33_4[49] <= 128'h01F00F80000000000000000000000000;
                                        char33_4[50] <= 128'h00F81F00000000000000000000000000;
                                        char33_4[51] <= 128'h007E7E00000000000000000000000000;
                                        char33_4[52] <= 128'h003FFC00000000000000000000000000;
                                        char33_4[53] <= 128'h000FF000000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//0
                                  4'd1: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h0000E000000000000000000000000000;
                                        char33_4[11] <= 128'h0001E000000000000000000000000000;
                                        char33_4[12] <= 128'h0003E000000000000000000000000000;
                                        char33_4[13] <= 128'h001FE000000000000000000000000000;
                                        char33_4[14] <= 128'h03FFE000000000000000000000000000;
                                        char33_4[15] <= 128'h03FFE000000000000000000000000000;
                                        char33_4[16] <= 128'h0007E000000000000000000000000000;
                                        char33_4[17] <= 128'h0007E000000000000000000000000000;
                                        char33_4[18] <= 128'h0007E000000000000000000000000000;
                                        char33_4[19] <= 128'h0007E000000000000000000000000000;
                                        char33_4[20] <= 128'h0007E000000000000000000000000000;
                                        char33_4[21] <= 128'h0007E000000000000000000000000000;
                                        char33_4[22] <= 128'h0007E000000000000000000000000000;
                                        char33_4[23] <= 128'h0007E000000000000000000000000000;
                                        char33_4[24] <= 128'h0007E000000000000000000000000000;
                                        char33_4[25] <= 128'h0007E000000000000000000000000000;
                                        char33_4[26] <= 128'h0007E000000000000000000000000000;
                                        char33_4[27] <= 128'h0007E000000000000000000000000000;
                                        char33_4[28] <= 128'h0007E000000000000000000000000000;
                                        char33_4[29] <= 128'h0007E000000000000000000000000000;
                                        char33_4[30] <= 128'h0007E000000000000000000000000000;
                                        char33_4[31] <= 128'h0007E000000000000000000000000000;
                                        char33_4[32] <= 128'h0007E000000000000000000000000000;
                                        char33_4[33] <= 128'h0007E000000000000000000000000000;
                                        char33_4[34] <= 128'h0007E000000000000000000000000000;
                                        char33_4[35] <= 128'h0007E000000000000000000000000000;
                                        char33_4[36] <= 128'h0007E000000000000000000000000000;
                                        char33_4[37] <= 128'h0007E000000000000000000000000000;
                                        char33_4[38] <= 128'h0007E000000000000000000000000000;
                                        char33_4[39] <= 128'h0007E000000000000000000000000000;
                                        char33_4[40] <= 128'h0007E000000000000000000000000000;
                                        char33_4[41] <= 128'h0007E000000000000000000000000000;
                                        char33_4[42] <= 128'h0007E000000000000000000000000000;
                                        char33_4[43] <= 128'h0007E000000000000000000000000000;
                                        char33_4[44] <= 128'h0007E000000000000000000000000000;
                                        char33_4[45] <= 128'h0007E000000000000000000000000000;
                                        char33_4[46] <= 128'h0007E000000000000000000000000000;
                                        char33_4[47] <= 128'h0007E000000000000000000000000000;
                                        char33_4[48] <= 128'h0007E000000000000000000000000000;
                                        char33_4[49] <= 128'h0007E000000000000000000000000000;
                                        char33_4[50] <= 128'h0007E000000000000000000000000000;
                                        char33_4[51] <= 128'h000FF800000000000000000000000000;
                                        char33_4[52] <= 128'h03FFFFC0000000000000000000000000;
                                        char33_4[53] <= 128'h03FFFFC0000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//1
                                  4'd2: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h001FFC00000000000000000000000000;
                                        char33_4[11] <= 128'h007FFF00000000000000000000000000;
                                        char33_4[12] <= 128'h01F83F80000000000000000000000000;
                                        char33_4[13] <= 128'h03E00FC0000000000000000000000000;
                                        char33_4[14] <= 128'h07C007E0000000000000000000000000;
                                        char33_4[15] <= 128'h078007E0000000000000000000000000;
                                        char33_4[16] <= 128'h0F8003F0000000000000000000000000;
                                        char33_4[17] <= 128'h0F8003F0000000000000000000000000;
                                        char33_4[18] <= 128'h1F8003F0000000000000000000000000;
                                        char33_4[19] <= 128'h1F8003F0000000000000000000000000;
                                        char33_4[20] <= 128'h1FC003F0000000000000000000000000;
                                        char33_4[21] <= 128'h1FC003F0000000000000000000000000;
                                        char33_4[22] <= 128'h1FC003F0000000000000000000000000;
                                        char33_4[23] <= 128'h0FC003F0000000000000000000000000;
                                        char33_4[24] <= 128'h07C003F0000000000000000000000000;
                                        char33_4[25] <= 128'h000003E0000000000000000000000000;
                                        char33_4[26] <= 128'h000007E0000000000000000000000000;
                                        char33_4[27] <= 128'h000007E0000000000000000000000000;
                                        char33_4[28] <= 128'h00000FC0000000000000000000000000;
                                        char33_4[29] <= 128'h00000F80000000000000000000000000;
                                        char33_4[30] <= 128'h00001F80000000000000000000000000;
                                        char33_4[31] <= 128'h00003F00000000000000000000000000;
                                        char33_4[32] <= 128'h00003E00000000000000000000000000;
                                        char33_4[33] <= 128'h00007C00000000000000000000000000;
                                        char33_4[34] <= 128'h0000F800000000000000000000000000;
                                        char33_4[35] <= 128'h0001F000000000000000000000000000;
                                        char33_4[36] <= 128'h0003E000000000000000000000000000;
                                        char33_4[37] <= 128'h0007C000000000000000000000000000;
                                        char33_4[38] <= 128'h000F8000000000000000000000000000;
                                        char33_4[39] <= 128'h001F0000000000000000000000000000;
                                        char33_4[40] <= 128'h003E0000000000000000000000000000;
                                        char33_4[41] <= 128'h007C0000000000000000000000000000;
                                        char33_4[42] <= 128'h00F80000000000000000000000000000;
                                        char33_4[43] <= 128'h01F00038000000000000000000000000;
                                        char33_4[44] <= 128'h01E00038000000000000000000000000;
                                        char33_4[45] <= 128'h03C00070000000000000000000000000;
                                        char33_4[46] <= 128'h07800070000000000000000000000000;
                                        char33_4[47] <= 128'h0F8000F0000000000000000000000000;
                                        char33_4[48] <= 128'h0F0000F0000000000000000000000000;
                                        char33_4[49] <= 128'h1E0003F0000000000000000000000000;
                                        char33_4[50] <= 128'h3FFFFFF0000000000000000000000000;
                                        char33_4[51] <= 128'h3FFFFFF0000000000000000000000000;
                                        char33_4[52] <= 128'h3FFFFFE0000000000000000000000000;
                                        char33_4[53] <= 128'h3FFFFFE0000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//2
                                  4'd3: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h003FF000000000000000000000000000;
                                        char33_4[11] <= 128'h00FFFC00000000000000000000000000;
                                        char33_4[12] <= 128'h01F07E00000000000000000000000000;
                                        char33_4[13] <= 128'h03C03F00000000000000000000000000;
                                        char33_4[14] <= 128'h07801F80000000000000000000000000;
                                        char33_4[15] <= 128'h0F800FC0000000000000000000000000;
                                        char33_4[16] <= 128'h0F800FC0000000000000000000000000;
                                        char33_4[17] <= 128'h0F8007E0000000000000000000000000;
                                        char33_4[18] <= 128'h0FC007E0000000000000000000000000;
                                        char33_4[19] <= 128'h0FC007E0000000000000000000000000;
                                        char33_4[20] <= 128'h0FC007E0000000000000000000000000;
                                        char33_4[21] <= 128'h07C007E0000000000000000000000000;
                                        char33_4[22] <= 128'h000007E0000000000000000000000000;
                                        char33_4[23] <= 128'h000007E0000000000000000000000000;
                                        char33_4[24] <= 128'h000007C0000000000000000000000000;
                                        char33_4[25] <= 128'h00000FC0000000000000000000000000;
                                        char33_4[26] <= 128'h00000F80000000000000000000000000;
                                        char33_4[27] <= 128'h00001F00000000000000000000000000;
                                        char33_4[28] <= 128'h00007E00000000000000000000000000;
                                        char33_4[29] <= 128'h0003FC00000000000000000000000000;
                                        char33_4[30] <= 128'h001FF000000000000000000000000000;
                                        char33_4[31] <= 128'h001FFC00000000000000000000000000;
                                        char33_4[32] <= 128'h0000FF00000000000000000000000000;
                                        char33_4[33] <= 128'h00001F80000000000000000000000000;
                                        char33_4[34] <= 128'h00000FC0000000000000000000000000;
                                        char33_4[35] <= 128'h000007E0000000000000000000000000;
                                        char33_4[36] <= 128'h000003E0000000000000000000000000;
                                        char33_4[37] <= 128'h000003F0000000000000000000000000;
                                        char33_4[38] <= 128'h000003F0000000000000000000000000;
                                        char33_4[39] <= 128'h000001F0000000000000000000000000;
                                        char33_4[40] <= 128'h000001F8000000000000000000000000;
                                        char33_4[41] <= 128'h000001F8000000000000000000000000;
                                        char33_4[42] <= 128'h078001F8000000000000000000000000;
                                        char33_4[43] <= 128'h0FC001F8000000000000000000000000;
                                        char33_4[44] <= 128'h1FC001F8000000000000000000000000;
                                        char33_4[45] <= 128'h1FC003F0000000000000000000000000;
                                        char33_4[46] <= 128'h1FC003F0000000000000000000000000;
                                        char33_4[47] <= 128'h1FC003E0000000000000000000000000;
                                        char33_4[48] <= 128'h0F8007E0000000000000000000000000;
                                        char33_4[49] <= 128'h0F8007C0000000000000000000000000;
                                        char33_4[50] <= 128'h07C01F80000000000000000000000000;
                                        char33_4[51] <= 128'h03F07F00000000000000000000000000;
                                        char33_4[52] <= 128'h01FFFE00000000000000000000000000;
                                        char33_4[53] <= 128'h003FF000000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//3
                                  4'd4: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h00001F00000000000000000000000000;
                                        char33_4[11] <= 128'h00001F00000000000000000000000000;
                                        char33_4[12] <= 128'h00003F00000000000000000000000000;
                                        char33_4[13] <= 128'h00003F00000000000000000000000000;
                                        char33_4[14] <= 128'h00007F00000000000000000000000000;
                                        char33_4[15] <= 128'h0000FF00000000000000000000000000;
                                        char33_4[16] <= 128'h0000FF00000000000000000000000000;
                                        char33_4[17] <= 128'h0001FF00000000000000000000000000;
                                        char33_4[18] <= 128'h0003FF00000000000000000000000000;
                                        char33_4[19] <= 128'h0003BF00000000000000000000000000;
                                        char33_4[20] <= 128'h0007BF00000000000000000000000000;
                                        char33_4[21] <= 128'h00073F00000000000000000000000000;
                                        char33_4[22] <= 128'h000F3F00000000000000000000000000;
                                        char33_4[23] <= 128'h001E3F00000000000000000000000000;
                                        char33_4[24] <= 128'h001C3F00000000000000000000000000;
                                        char33_4[25] <= 128'h003C3F00000000000000000000000000;
                                        char33_4[26] <= 128'h00783F00000000000000000000000000;
                                        char33_4[27] <= 128'h00783F00000000000000000000000000;
                                        char33_4[28] <= 128'h00F03F00000000000000000000000000;
                                        char33_4[29] <= 128'h00E03F00000000000000000000000000;
                                        char33_4[30] <= 128'h01E03F00000000000000000000000000;
                                        char33_4[31] <= 128'h03C03F00000000000000000000000000;
                                        char33_4[32] <= 128'h03803F00000000000000000000000000;
                                        char33_4[33] <= 128'h07803F00000000000000000000000000;
                                        char33_4[34] <= 128'h0F003F00000000000000000000000000;
                                        char33_4[35] <= 128'h0F003F00000000000000000000000000;
                                        char33_4[36] <= 128'h1E003F00000000000000000000000000;
                                        char33_4[37] <= 128'h1C003F00000000000000000000000000;
                                        char33_4[38] <= 128'h3C003F00000000000000000000000000;
                                        char33_4[39] <= 128'h7FFFFFFE000000000000000000000000;
                                        char33_4[40] <= 128'h7FFFFFFE000000000000000000000000;
                                        char33_4[41] <= 128'h00003F00000000000000000000000000;
                                        char33_4[42] <= 128'h00003F00000000000000000000000000;
                                        char33_4[43] <= 128'h00003F00000000000000000000000000;
                                        char33_4[44] <= 128'h00003F00000000000000000000000000;
                                        char33_4[45] <= 128'h00003F00000000000000000000000000;
                                        char33_4[46] <= 128'h00003F00000000000000000000000000;
                                        char33_4[47] <= 128'h00003F00000000000000000000000000;
                                        char33_4[48] <= 128'h00003F00000000000000000000000000;
                                        char33_4[49] <= 128'h00003F00000000000000000000000000;
                                        char33_4[50] <= 128'h00003F00000000000000000000000000;
                                        char33_4[51] <= 128'h00007F80000000000000000000000000;
                                        char33_4[52] <= 128'h000FFFFC000000000000000000000000;
                                        char33_4[53] <= 128'h000FFFFC000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//4
                                  4'd5: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h00000000000000000000000000000000;
                                        char33_4[11] <= 128'h03FFFFF0000000000000000000000000;
                                        char33_4[12] <= 128'h03FFFFF0000000000000000000000000;
                                        char33_4[13] <= 128'h03FFFFF0000000000000000000000000;
                                        char33_4[14] <= 128'h03FFFFE0000000000000000000000000;
                                        char33_4[15] <= 128'h03800000000000000000000000000000;
                                        char33_4[16] <= 128'h03800000000000000000000000000000;
                                        char33_4[17] <= 128'h03800000000000000000000000000000;
                                        char33_4[18] <= 128'h03800000000000000000000000000000;
                                        char33_4[19] <= 128'h03800000000000000000000000000000;
                                        char33_4[20] <= 128'h07800000000000000000000000000000;
                                        char33_4[21] <= 128'h07800000000000000000000000000000;
                                        char33_4[22] <= 128'h07800000000000000000000000000000;
                                        char33_4[23] <= 128'h07800000000000000000000000000000;
                                        char33_4[24] <= 128'h07800000000000000000000000000000;
                                        char33_4[25] <= 128'h07800000000000000000000000000000;
                                        char33_4[26] <= 128'h078FF800000000000000000000000000;
                                        char33_4[27] <= 128'h073FFE00000000000000000000000000;
                                        char33_4[28] <= 128'h077FFF80000000000000000000000000;
                                        char33_4[29] <= 128'h07FC3F80000000000000000000000000;
                                        char33_4[30] <= 128'h07E00FC0000000000000000000000000;
                                        char33_4[31] <= 128'h07C007E0000000000000000000000000;
                                        char33_4[32] <= 128'h078007E0000000000000000000000000;
                                        char33_4[33] <= 128'h078003F0000000000000000000000000;
                                        char33_4[34] <= 128'h000003F0000000000000000000000000;
                                        char33_4[35] <= 128'h000001F0000000000000000000000000;
                                        char33_4[36] <= 128'h000001F8000000000000000000000000;
                                        char33_4[37] <= 128'h000001F8000000000000000000000000;
                                        char33_4[38] <= 128'h000001F8000000000000000000000000;
                                        char33_4[39] <= 128'h000001F8000000000000000000000000;
                                        char33_4[40] <= 128'h000001F8000000000000000000000000;
                                        char33_4[41] <= 128'h078001F8000000000000000000000000;
                                        char33_4[42] <= 128'h0FC001F8000000000000000000000000;
                                        char33_4[43] <= 128'h1FC001F0000000000000000000000000;
                                        char33_4[44] <= 128'h1FC001F0000000000000000000000000;
                                        char33_4[45] <= 128'h1FC003F0000000000000000000000000;
                                        char33_4[46] <= 128'h1F8003F0000000000000000000000000;
                                        char33_4[47] <= 128'h1F8003E0000000000000000000000000;
                                        char33_4[48] <= 128'h0F8007E0000000000000000000000000;
                                        char33_4[49] <= 128'h078007C0000000000000000000000000;
                                        char33_4[50] <= 128'h07C01F80000000000000000000000000;
                                        char33_4[51] <= 128'h03F83F00000000000000000000000000;
                                        char33_4[52] <= 128'h00FFFE00000000000000000000000000;
                                        char33_4[53] <= 128'h003FF800000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//5
                                  4'd6: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h0007FE00000000000000000000000000;
                                        char33_4[11] <= 128'h001FFF80000000000000000000000000;
                                        char33_4[12] <= 128'h003F0FC0000000000000000000000000;
                                        char33_4[13] <= 128'h007C07C0000000000000000000000000;
                                        char33_4[14] <= 128'h00F807E0000000000000000000000000;
                                        char33_4[15] <= 128'h01F007E0000000000000000000000000;
                                        char33_4[16] <= 128'h03E007E0000000000000000000000000;
                                        char33_4[17] <= 128'h03C007E0000000000000000000000000;
                                        char33_4[18] <= 128'h07C003C0000000000000000000000000;
                                        char33_4[19] <= 128'h07C00000000000000000000000000000;
                                        char33_4[20] <= 128'h0FC00000000000000000000000000000;
                                        char33_4[21] <= 128'h0F800000000000000000000000000000;
                                        char33_4[22] <= 128'h0F800000000000000000000000000000;
                                        char33_4[23] <= 128'h1F800000000000000000000000000000;
                                        char33_4[24] <= 128'h1F800000000000000000000000000000;
                                        char33_4[25] <= 128'h1F800000000000000000000000000000;
                                        char33_4[26] <= 128'h1F87FE00000000000000000000000000;
                                        char33_4[27] <= 128'h1F9FFF80000000000000000000000000;
                                        char33_4[28] <= 128'h1FBFFFC0000000000000000000000000;
                                        char33_4[29] <= 128'h3FFE1FC0000000000000000000000000;
                                        char33_4[30] <= 128'h3FF807E0000000000000000000000000;
                                        char33_4[31] <= 128'h3FE003F0000000000000000000000000;
                                        char33_4[32] <= 128'h3FE003F0000000000000000000000000;
                                        char33_4[33] <= 128'h3FC001F8000000000000000000000000;
                                        char33_4[34] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[35] <= 128'h3F8001F8000000000000000000000000;
                                        char33_4[36] <= 128'h3F8000F8000000000000000000000000;
                                        char33_4[37] <= 128'h3F8000F8000000000000000000000000;
                                        char33_4[38] <= 128'h3F8000F8000000000000000000000000;
                                        char33_4[39] <= 128'h1F8000F8000000000000000000000000;
                                        char33_4[40] <= 128'h1F8000F8000000000000000000000000;
                                        char33_4[41] <= 128'h1F8000F8000000000000000000000000;
                                        char33_4[42] <= 128'h1F8000F8000000000000000000000000;
                                        char33_4[43] <= 128'h1F8000F8000000000000000000000000;
                                        char33_4[44] <= 128'h0FC001F8000000000000000000000000;
                                        char33_4[45] <= 128'h0FC001F8000000000000000000000000;
                                        char33_4[46] <= 128'h0FC001F0000000000000000000000000;
                                        char33_4[47] <= 128'h07E001F0000000000000000000000000;
                                        char33_4[48] <= 128'h03E003E0000000000000000000000000;
                                        char33_4[49] <= 128'h03F003E0000000000000000000000000;
                                        char33_4[50] <= 128'h01F807C0000000000000000000000000;
                                        char33_4[51] <= 128'h00FE1F80000000000000000000000000;
                                        char33_4[52] <= 128'h007FFE00000000000000000000000000;
                                        char33_4[53] <= 128'h001FF800000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//6
                                  4'd7: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h00000000000000000000000000000000;
                                        char33_4[11] <= 128'h07FFFFF8000000000000000000000000;
                                        char33_4[12] <= 128'h07FFFFF8000000000000000000000000;
                                        char33_4[13] <= 128'h07FFFFF8000000000000000000000000;
                                        char33_4[14] <= 128'h0FFFFFF0000000000000000000000000;
                                        char33_4[15] <= 128'h0FC000E0000000000000000000000000;
                                        char33_4[16] <= 128'h0F8001E0000000000000000000000000;
                                        char33_4[17] <= 128'h0F0001C0000000000000000000000000;
                                        char33_4[18] <= 128'h0E0003C0000000000000000000000000;
                                        char33_4[19] <= 128'h0E000780000000000000000000000000;
                                        char33_4[20] <= 128'h1E000780000000000000000000000000;
                                        char33_4[21] <= 128'h1C000F00000000000000000000000000;
                                        char33_4[22] <= 128'h00000F00000000000000000000000000;
                                        char33_4[23] <= 128'h00001E00000000000000000000000000;
                                        char33_4[24] <= 128'h00001E00000000000000000000000000;
                                        char33_4[25] <= 128'h00003C00000000000000000000000000;
                                        char33_4[26] <= 128'h00003C00000000000000000000000000;
                                        char33_4[27] <= 128'h00007800000000000000000000000000;
                                        char33_4[28] <= 128'h00007800000000000000000000000000;
                                        char33_4[29] <= 128'h0000F800000000000000000000000000;
                                        char33_4[30] <= 128'h0000F000000000000000000000000000;
                                        char33_4[31] <= 128'h0001F000000000000000000000000000;
                                        char33_4[32] <= 128'h0001E000000000000000000000000000;
                                        char33_4[33] <= 128'h0003E000000000000000000000000000;
                                        char33_4[34] <= 128'h0003E000000000000000000000000000;
                                        char33_4[35] <= 128'h0003E000000000000000000000000000;
                                        char33_4[36] <= 128'h0007C000000000000000000000000000;
                                        char33_4[37] <= 128'h0007C000000000000000000000000000;
                                        char33_4[38] <= 128'h0007C000000000000000000000000000;
                                        char33_4[39] <= 128'h000FC000000000000000000000000000;
                                        char33_4[40] <= 128'h000FC000000000000000000000000000;
                                        char33_4[41] <= 128'h000FC000000000000000000000000000;
                                        char33_4[42] <= 128'h000FC000000000000000000000000000;
                                        char33_4[43] <= 128'h001FC000000000000000000000000000;
                                        char33_4[44] <= 128'h001FC000000000000000000000000000;
                                        char33_4[45] <= 128'h001FC000000000000000000000000000;
                                        char33_4[46] <= 128'h001FC000000000000000000000000000;
                                        char33_4[47] <= 128'h001FC000000000000000000000000000;
                                        char33_4[48] <= 128'h001FC000000000000000000000000000;
                                        char33_4[49] <= 128'h001FC000000000000000000000000000;
                                        char33_4[50] <= 128'h001FC000000000000000000000000000;
                                        char33_4[51] <= 128'h001FC000000000000000000000000000;
                                        char33_4[52] <= 128'h001FC000000000000000000000000000;
                                        char33_4[53] <= 128'h000F8000000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//7
                                  4'd8: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h003FF800000000000000000000000000;
                                        char33_4[11] <= 128'h00FFFE00000000000000000000000000;
                                        char33_4[12] <= 128'h01F81F80000000000000000000000000;
                                        char33_4[13] <= 128'h03E00FC0000000000000000000000000;
                                        char33_4[14] <= 128'h07C003E0000000000000000000000000;
                                        char33_4[15] <= 128'h0F8003E0000000000000000000000000;
                                        char33_4[16] <= 128'h0F8001F0000000000000000000000000;
                                        char33_4[17] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[18] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[19] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[20] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[21] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[22] <= 128'h1F8001F0000000000000000000000000;
                                        char33_4[23] <= 128'h1FC001F0000000000000000000000000;
                                        char33_4[24] <= 128'h0FC001F0000000000000000000000000;
                                        char33_4[25] <= 128'h0FF003E0000000000000000000000000;
                                        char33_4[26] <= 128'h07F803C0000000000000000000000000;
                                        char33_4[27] <= 128'h03FE0F80000000000000000000000000;
                                        char33_4[28] <= 128'h01FF9F00000000000000000000000000;
                                        char33_4[29] <= 128'h00FFFE00000000000000000000000000;
                                        char33_4[30] <= 128'h003FF800000000000000000000000000;
                                        char33_4[31] <= 128'h007FFC00000000000000000000000000;
                                        char33_4[32] <= 128'h01F7FF00000000000000000000000000;
                                        char33_4[33] <= 128'h03E1FF80000000000000000000000000;
                                        char33_4[34] <= 128'h07C07FC0000000000000000000000000;
                                        char33_4[35] <= 128'h0F801FE0000000000000000000000000;
                                        char33_4[36] <= 128'h0F800FE0000000000000000000000000;
                                        char33_4[37] <= 128'h1F0007F0000000000000000000000000;
                                        char33_4[38] <= 128'h1F0003F0000000000000000000000000;
                                        char33_4[39] <= 128'h3E0001F8000000000000000000000000;
                                        char33_4[40] <= 128'h3E0001F8000000000000000000000000;
                                        char33_4[41] <= 128'h3E0001F8000000000000000000000000;
                                        char33_4[42] <= 128'h3E0000F8000000000000000000000000;
                                        char33_4[43] <= 128'h3E0000F8000000000000000000000000;
                                        char33_4[44] <= 128'h3E0000F8000000000000000000000000;
                                        char33_4[45] <= 128'h3E0000F8000000000000000000000000;
                                        char33_4[46] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[47] <= 128'h1F0001F0000000000000000000000000;
                                        char33_4[48] <= 128'h0F8003E0000000000000000000000000;
                                        char33_4[49] <= 128'h0FC003E0000000000000000000000000;
                                        char33_4[50] <= 128'h07E007C0000000000000000000000000;
                                        char33_4[51] <= 128'h01F83F80000000000000000000000000;
                                        char33_4[52] <= 128'h00FFFE00000000000000000000000000;
                                        char33_4[53] <= 128'h003FF800000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//8
                                  4'd9: begin
                                        char33_4[0] <= 128'h00000000000000000000000000000000;
                                        char33_4[1] <= 128'h00000000000000000000000000000000;
                                        char33_4[2] <= 128'h00000000000000000000000000000000;
                                        char33_4[3] <= 128'h00000000000000000000000000000000;
                                        char33_4[4] <= 128'h00000000000000000000000000000000;
                                        char33_4[5] <= 128'h00000000000000000000000000000000;
                                        char33_4[6] <= 128'h00000000000000000000000000000000;
                                        char33_4[7] <= 128'h00000000000000000000000000000000;
                                        char33_4[8] <= 128'h00000000000000000000000000000000;
                                        char33_4[9] <= 128'h00000000000000000000000000000000;
                                        char33_4[10] <= 128'h003FF000000000000000000000000000;
                                        char33_4[11] <= 128'h00FFFC00000000000000000000000000;
                                        char33_4[12] <= 128'h01F83F00000000000000000000000000;
                                        char33_4[13] <= 128'h03E01F80000000000000000000000000;
                                        char33_4[14] <= 128'h07C00F80000000000000000000000000;
                                        char33_4[15] <= 128'h0FC007C0000000000000000000000000;
                                        char33_4[16] <= 128'h0F8003E0000000000000000000000000;
                                        char33_4[17] <= 128'h1F8003E0000000000000000000000000;
                                        char33_4[18] <= 128'h1F0003F0000000000000000000000000;
                                        char33_4[19] <= 128'h1F0003F0000000000000000000000000;
                                        char33_4[20] <= 128'h3F0001F0000000000000000000000000;
                                        char33_4[21] <= 128'h3F0001F0000000000000000000000000;
                                        char33_4[22] <= 128'h3F0001F8000000000000000000000000;
                                        char33_4[23] <= 128'h3F0001F8000000000000000000000000;
                                        char33_4[24] <= 128'h3F0001F8000000000000000000000000;
                                        char33_4[25] <= 128'h3F0001F8000000000000000000000000;
                                        char33_4[26] <= 128'h3F0001F8000000000000000000000000;
                                        char33_4[27] <= 128'h3F0001F8000000000000000000000000;
                                        char33_4[28] <= 128'h3F0003F8000000000000000000000000;
                                        char33_4[29] <= 128'h1F8003F8000000000000000000000000;
                                        char33_4[30] <= 128'h1F8007F8000000000000000000000000;
                                        char33_4[31] <= 128'h1F800FF8000000000000000000000000;
                                        char33_4[32] <= 128'h0FC01FF8000000000000000000000000;
                                        char33_4[33] <= 128'h0FE03FF8000000000000000000000000;
                                        char33_4[34] <= 128'h07F8FDF8000000000000000000000000;
                                        char33_4[35] <= 128'h03FFF9F8000000000000000000000000;
                                        char33_4[36] <= 128'h01FFF1F8000000000000000000000000;
                                        char33_4[37] <= 128'h003F83F8000000000000000000000000;
                                        char33_4[38] <= 128'h000003F0000000000000000000000000;
                                        char33_4[39] <= 128'h000003F0000000000000000000000000;
                                        char33_4[40] <= 128'h000003F0000000000000000000000000;
                                        char33_4[41] <= 128'h000003F0000000000000000000000000;
                                        char33_4[42] <= 128'h000007E0000000000000000000000000;
                                        char33_4[43] <= 128'h000007E0000000000000000000000000;
                                        char33_4[44] <= 128'h000007C0000000000000000000000000;
                                        char33_4[45] <= 128'h03C007C0000000000000000000000000;
                                        char33_4[46] <= 128'h07C00F80000000000000000000000000;
                                        char33_4[47] <= 128'h0FE00F80000000000000000000000000;
                                        char33_4[48] <= 128'h0FE01F00000000000000000000000000;
                                        char33_4[49] <= 128'h0FE03E00000000000000000000000000;
                                        char33_4[50] <= 128'h07E07E00000000000000000000000000;
                                        char33_4[51] <= 128'h07F1F800000000000000000000000000;
                                        char33_4[52] <= 128'h03FFF000000000000000000000000000;
                                        char33_4[53] <= 128'h00FFC000000000000000000000000000;
                                        char33_4[54] <= 128'h00000000000000000000000000000000;
                                        char33_4[55] <= 128'h00000000000000000000000000000000;
                                        char33_4[56] <= 128'h00000000000000000000000000000000;
                                        char33_4[57] <= 128'h00000000000000000000000000000000;
                                        char33_4[58] <= 128'h00000000000000000000000000000000;
                                        char33_4[59] <= 128'h00000000000000000000000000000000;
                                        char33_4[60] <= 128'h00000000000000000000000000000000;
                                        char33_4[61] <= 128'h00000000000000000000000000000000;
                                        char33_4[62] <= 128'h00000000000000000000000000000000;
                                        char33_4[63] <= 128'h00000000000000000000000000000000;
                                  end//9
                                  default: begin
                                      char33_4[0] <= char33_4[0];
                                      char33_4[1] <= char33_4[1];
                                      char33_4[2] <= char33_4[2];
                                      char33_4[3] <= char33_4[3];
                                      char33_4[4] <= char33_4[4];
                                      char33_4[5] <= char33_4[5];
                                      char33_4[6] <= char33_4[6];
                                      char33_4[7] <= char33_4[7];
                                      char33_4[8] <= char33_4[8];
                                      char33_4[9] <= char33_4[9];
                                      char33_4[10] <= char33_4[10];
                                      char33_4[11] <= char33_4[11];
                                      char33_4[12] <= char33_4[12];
                                      char33_4[13] <= char33_4[13];
                                      char33_4[14] <= char33_4[14];
                                      char33_4[15] <= char33_4[15];
                                      char33_4[16] <= char33_4[16];
                                      char33_4[17] <= char33_4[17];
                                      char33_4[18] <= char33_4[18];
                                      char33_4[19] <= char33_4[19];
                                      char33_4[20] <= char33_4[20];
                                      char33_4[21] <= char33_4[21];
                                      char33_4[22] <= char33_4[22];
                                      char33_4[23] <= char33_4[23];
                                      char33_4[24] <= char33_4[24];
                                      char33_4[25] <= char33_4[25];
                                      char33_4[26] <= char33_4[26];
                                      char33_4[27] <= char33_4[27];
                                      char33_4[28] <= char33_4[28];
                                      char33_4[29] <= char33_4[29];
                                      char33_4[30] <= char33_4[30];
                                      char33_4[31] <= char33_4[31];
                                      char33_4[32] <= char33_4[32];
                                      char33_4[33] <= char33_4[33];
                                      char33_4[34] <= char33_4[34];
                                      char33_4[35] <= char33_4[35];
                                      char33_4[36] <= char33_4[36];
                                      char33_4[37] <= char33_4[37];
                                      char33_4[38] <= char33_4[38];
                                      char33_4[39] <= char33_4[39];
                                      char33_4[40] <= char33_4[40];
                                      char33_4[41] <= char33_4[41];
                                      char33_4[42] <= char33_4[42];
                                      char33_4[43] <= char33_4[43];
                                      char33_4[44] <= char33_4[44];
                                      char33_4[45] <= char33_4[45];
                                      char33_4[46] <= char33_4[46];
                                      char33_4[47] <= char33_4[47];
                                      char33_4[48] <= char33_4[48];
                                      char33_4[49] <= char33_4[49];
                                      char33_4[50] <= char33_4[50];
                                      char33_4[51] <= char33_4[51];
                                      char33_4[52] <= char33_4[52];
                                      char33_4[53] <= char33_4[53];
                                      char33_4[54] <= char33_4[54];
                                      char33_4[55] <= char33_4[55];
                                      char33_4[56] <= char33_4[56];
                                      char33_4[57] <= char33_4[57];
                                      char33_4[58] <= char33_4[58];
                                      char33_4[59] <= char33_4[59];
                                      char33_4[60] <= char33_4[60];
                                      char33_4[61] <= char33_4[61];
                                      char33_4[62] <= char33_4[62];
                                      char33_4[63] <= char33_4[63];
                                  end
                              endcase
                      
         case(a2/w1)
                                  4'd0: begin
                                      char44_0[  0] <= 32'h00000000;
                                      char44_0[  1] <= 32'h00000000;
                                      char44_0[  2] <= 32'h00000000;
                                      char44_0[  3] <= 32'h00000000;
                                      char44_0[  4] <= 32'h00000000;
                                      char44_0[  5] <= 32'h00000000;
                                      char44_0[  6] <= 32'h00000000;
                                      char44_0[  7] <= 32'h00000000;
                                      char44_0[  8] <= 32'h00000000;
                                      char44_0[  9] <= 32'h00000000;
                                      char44_0[10] <= 32'h000FF000;
                                      char44_0[11] <= 32'h003FFC00;
                                      char44_0[12] <= 32'h007E7E00;
                                      char44_0[13] <= 32'h00F81F00;
                                      char44_0[14] <= 32'h01F00F80;
                                      char44_0[15] <= 32'h03F00FC0;
                                      char44_0[16] <= 32'h03E007C0;
                                      char44_0[17] <= 32'h07E007E0;
                                      char44_0[18] <= 32'h07C003E0;
                                      char44_0[19] <= 32'h0FC003F0;
                                      char44_0[20] <= 32'h0FC003F0;
                                      char44_0[21] <= 32'h0FC003F0;
                                      char44_0[22] <= 32'h1F8001F8;
                                      char44_0[23] <= 32'h1F8001F8;
                                      char44_0[24] <= 32'h1F8001F8;
                                      char44_0[25] <= 32'h1F8001F8;
                                      char44_0[26] <= 32'h1F8001F8;
                                      char44_0[27] <= 32'h3F8001F8;
                                      char44_0[28] <= 32'h3F8001F8;
                                      char44_0[29] <= 32'h3F8001F8;
                                      char44_0[30] <= 32'h3F8001F8;
                                      char44_0[31] <= 32'h3F8001F8;
                                      char44_0[32] <= 32'h3F8001F8;
                                      char44_0[33] <= 32'h3F8001F8;
                                      char44_0[34] <= 32'h3F8001F8;
                                      char44_0[35] <= 32'h3F8001F8;
                                      char44_0[36] <= 32'h3F8001F8;
                                      char44_0[37] <= 32'h1F8001F8;
                                      char44_0[38] <= 32'h1F8001F8;
                                      char44_0[39] <= 32'h1F8001F8;
                                      char44_0[40] <= 32'h1F8001F8;
                                      char44_0[41] <= 32'h1F8001F0;
                                      char44_0[42] <= 32'h0F8003F0;
                                      char44_0[43] <= 32'h0FC003F0;
                                      char44_0[44] <= 32'h0FC003F0;
                                      char44_0[45] <= 32'h07C003E0;
                                      char44_0[46] <= 32'h07E007E0;
                                      char44_0[47] <= 32'h03E007C0;
                                      char44_0[48] <= 32'h03F00FC0;
                                      char44_0[49] <= 32'h01F00F80;
                                      char44_0[50] <= 32'h00F81F00;
                                      char44_0[51] <= 32'h007E7E00;
                                      char44_0[52] <= 32'h003FFC00;
                                      char44_0[53] <= 32'h000FF000;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//0
                                  4'd1: begin
                                      char44_0[  0] <= 32'h00000000;
                                      char44_0[  1] <= 32'h00000000;
                                      char44_0[  2] <= 32'h00000000;
                                      char44_0[  3] <= 32'h00000000;
                                      char44_0[  4] <= 32'h00000000;
                                      char44_0[  5] <= 32'h00000000;
                                      char44_0[  6] <= 32'h00000000;
                                      char44_0[  7] <= 32'h00000000;
                                      char44_0[  8] <= 32'h00000000;
                                      char44_0[  9] <= 32'h00000000;
                                      char44_0[10] <= 32'h0000E000;
                                      char44_0[11] <= 32'h0001E000;
                                      char44_0[12] <= 32'h0003E000;
                                      char44_0[13] <= 32'h001FE000;
                                      char44_0[14] <= 32'h03FFE000;
                                      char44_0[15] <= 32'h03FFE000;
                                      char44_0[16] <= 32'h0007E000;
                                      char44_0[17] <= 32'h0007E000;
                                      char44_0[18] <= 32'h0007E000;
                                      char44_0[19] <= 32'h0007E000;
                                      char44_0[20] <= 32'h0007E000;
                                      char44_0[21] <= 32'h0007E000;
                                      char44_0[22] <= 32'h0007E000;
                                      char44_0[23] <= 32'h0007E000;
                                      char44_0[24] <= 32'h0007E000;
                                      char44_0[25] <= 32'h0007E000;
                                      char44_0[26] <= 32'h0007E000;
                                      char44_0[27] <= 32'h0007E000;
                                      char44_0[28] <= 32'h0007E000;
                                      char44_0[29] <= 32'h0007E000;
                                      char44_0[30] <= 32'h0007E000;
                                      char44_0[31] <= 32'h0007E000;
                                      char44_0[32] <= 32'h0007E000;
                                      char44_0[33] <= 32'h0007E000;
                                      char44_0[34] <= 32'h0007E000;
                                      char44_0[35] <= 32'h0007E000;
                                      char44_0[36] <= 32'h0007E000;
                                      char44_0[37] <= 32'h0007E000;
                                      char44_0[38] <= 32'h0007E000;
                                      char44_0[39] <= 32'h0007E000;
                                      char44_0[40] <= 32'h0007E000;
                                      char44_0[41] <= 32'h0007E000;
                                      char44_0[42] <= 32'h0007E000;
                                      char44_0[43] <= 32'h0007E000;
                                      char44_0[44] <= 32'h0007E000;
                                      char44_0[45] <= 32'h0007E000;
                                      char44_0[46] <= 32'h0007E000;
                                      char44_0[47] <= 32'h0007E000;
                                      char44_0[48] <= 32'h0007E000;
                                      char44_0[49] <= 32'h0007E000;
                                      char44_0[50] <= 32'h0007E000;
                                      char44_0[51] <= 32'h000FF800;
                                      char44_0[52] <= 32'h03FFFFC0;
                                      char44_0[53] <= 32'h03FFFFC0;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//1
                                  4'd2: begin
                                      char44_0[  0] <= 32'h00000000;
                                      char44_0[  1] <= 32'h00000000;
                                      char44_0[  2] <= 32'h00000000;
                                      char44_0[  3] <= 32'h00000000;
                                      char44_0[  4] <= 32'h00000000;
                                      char44_0[  5] <= 32'h00000000;
                                      char44_0[  6] <= 32'h00000000;
                                      char44_0[  7] <= 32'h00000000;
                                      char44_0[  8] <= 32'h00000000;
                                      char44_0[  9] <= 32'h00000000;
                                      char44_0[10] <= 32'h001FFC00;
                                      char44_0[11] <= 32'h007FFF00;
                                      char44_0[12] <= 32'h01F83F80;
                                      char44_0[13] <= 32'h03E00FC0;
                                      char44_0[14] <= 32'h07C007E0;
                                      char44_0[15] <= 32'h078007E0;
                                      char44_0[16] <= 32'h0F8003F0;
                                      char44_0[17] <= 32'h0F8003F0;
                                      char44_0[18] <= 32'h1F8003F0;
                                      char44_0[19] <= 32'h1F8003F0;
                                      char44_0[20] <= 32'h1FC003F0;
                                      char44_0[21] <= 32'h1FC003F0;
                                      char44_0[22] <= 32'h1FC003F0;
                                      char44_0[23] <= 32'h0FC003F0;
                                      char44_0[24] <= 32'h07C003F0;
                                      char44_0[25] <= 32'h000003E0;
                                      char44_0[26] <= 32'h000007E0;
                                      char44_0[27] <= 32'h000007E0;
                                      char44_0[28] <= 32'h00000FC0;
                                      char44_0[29] <= 32'h00000F80;
                                      char44_0[30] <= 32'h00001F80;
                                      char44_0[31] <= 32'h00003F00;
                                      char44_0[32] <= 32'h00003E00;
                                      char44_0[33] <= 32'h00007C00;
                                      char44_0[34] <= 32'h0000F800;
                                      char44_0[35] <= 32'h0001F000;
                                      char44_0[36] <= 32'h0003E000;
                                      char44_0[37] <= 32'h0007C000;
                                      char44_0[38] <= 32'h000F8000;
                                      char44_0[39] <= 32'h001F0000;
                                      char44_0[40] <= 32'h003E0000;
                                      char44_0[41] <= 32'h007C0000;
                                      char44_0[42] <= 32'h00F80000;
                                      char44_0[43] <= 32'h01F00038;
                                      char44_0[44] <= 32'h01E00038;
                                      char44_0[45] <= 32'h03C00070;
                                      char44_0[46] <= 32'h07800070;
                                      char44_0[47] <= 32'h0F8000F0;
                                      char44_0[48] <= 32'h0F0000F0;
                                      char44_0[49] <= 32'h1E0003F0;
                                      char44_0[50] <= 32'h3FFFFFF0;
                                      char44_0[51] <= 32'h3FFFFFF0;
                                      char44_0[52] <= 32'h3FFFFFE0;
                                      char44_0[53] <= 32'h3FFFFFE0;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//2
                                  4'd3: begin
                                      char44_0[  0] <= 32'h00000000;
                                      char44_0[  1] <= 32'h00000000;
                                      char44_0[  2] <= 32'h00000000;
                                      char44_0[  3] <= 32'h00000000;
                                      char44_0[  4] <= 32'h00000000;
                                      char44_0[  5] <= 32'h00000000;
                                      char44_0[  6] <= 32'h00000000;
                                      char44_0[  7] <= 32'h00000000;
                                      char44_0[  8] <= 32'h00000000;
                                      char44_0[  9] <= 32'h00000000;
                                      char44_0[10] <= 32'h003FF000;
                                      char44_0[11] <= 32'h00FFFC00;
                                      char44_0[12] <= 32'h01F07E00;
                                      char44_0[13] <= 32'h03C03F00;
                                      char44_0[14] <= 32'h07801F80;
                                      char44_0[15] <= 32'h0F800FC0;
                                      char44_0[16] <= 32'h0F800FC0;
                                      char44_0[17] <= 32'h0F8007E0;
                                      char44_0[18] <= 32'h0FC007E0;
                                      char44_0[19] <= 32'h0FC007E0;
                                      char44_0[20] <= 32'h0FC007E0;
                                      char44_0[21] <= 32'h07C007E0;
                                      char44_0[22] <= 32'h000007E0;
                                      char44_0[23] <= 32'h000007E0;
                                      char44_0[24] <= 32'h000007C0;
                                      char44_0[25] <= 32'h00000FC0;
                                      char44_0[26] <= 32'h00000F80;
                                      char44_0[27] <= 32'h00001F00;
                                      char44_0[28] <= 32'h00007E00;
                                      char44_0[29] <= 32'h0003FC00;
                                      char44_0[30] <= 32'h001FF000;
                                      char44_0[31] <= 32'h001FFC00;
                                      char44_0[32] <= 32'h0000FF00;
                                      char44_0[33] <= 32'h00001F80;
                                      char44_0[34] <= 32'h00000FC0;
                                      char44_0[35] <= 32'h000007E0;
                                      char44_0[36] <= 32'h000003E0;
                                      char44_0[37] <= 32'h000003F0;
                                      char44_0[38] <= 32'h000003F0;
                                      char44_0[39] <= 32'h000001F0;
                                      char44_0[40] <= 32'h000001F8;
                                      char44_0[41] <= 32'h000001F8;
                                      char44_0[42] <= 32'h078001F8;
                                      char44_0[43] <= 32'h0FC001F8;
                                      char44_0[44] <= 32'h1FC001F8;
                                      char44_0[45] <= 32'h1FC003F0;
                                      char44_0[46] <= 32'h1FC003F0;
                                      char44_0[47] <= 32'h1FC003E0;
                                      char44_0[48] <= 32'h0F8007E0;
                                      char44_0[49] <= 32'h0F8007C0;
                                      char44_0[50] <= 32'h07C01F80;
                                      char44_0[51] <= 32'h03F07F00;
                                      char44_0[52] <= 32'h01FFFE00;
                                      char44_0[53] <= 32'h003FF000;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//3
                                  4'd4: begin
                                      char44_0[  0] <= 32'h00000000;
                                      char44_0[  1] <= 32'h00000000;
                                      char44_0[  2] <= 32'h00000000;
                                      char44_0[  3] <= 32'h00000000;
                                      char44_0[  4] <= 32'h00000000;
                                      char44_0[  5] <= 32'h00000000;
                                      char44_0[  6] <= 32'h00000000;
                                      char44_0[  7] <= 32'h00000000;
                                      char44_0[  8] <= 32'h00000000;
                                      char44_0[  9] <= 32'h00000000;
                                      char44_0[10] <= 32'h00001F00;
                                      char44_0[11] <= 32'h00001F00;
                                      char44_0[12] <= 32'h00003F00;
                                      char44_0[13] <= 32'h00003F00;
                                      char44_0[14] <= 32'h00007F00;
                                      char44_0[15] <= 32'h0000FF00;
                                      char44_0[16] <= 32'h0000FF00;
                                      char44_0[17] <= 32'h0001FF00;
                                      char44_0[18] <= 32'h0003FF00;
                                      char44_0[19] <= 32'h0003BF00;
                                      char44_0[20] <= 32'h0007BF00;
                                      char44_0[21] <= 32'h00073F00;
                                      char44_0[22] <= 32'h000F3F00;
                                      char44_0[23] <= 32'h001E3F00;
                                      char44_0[24] <= 32'h001C3F00;
                                      char44_0[25] <= 32'h003C3F00;
                                      char44_0[26] <= 32'h00783F00;
                                      char44_0[27] <= 32'h00783F00;
                                      char44_0[28] <= 32'h00F03F00;
                                      char44_0[29] <= 32'h00E03F00;
                                      char44_0[30] <= 32'h01E03F00;
                                      char44_0[31] <= 32'h03C03F00;
                                      char44_0[32] <= 32'h03803F00;
                                      char44_0[33] <= 32'h07803F00;
                                      char44_0[34] <= 32'h0F003F00;
                                      char44_0[35] <= 32'h0F003F00;
                                      char44_0[36] <= 32'h1E003F00;
                                      char44_0[37] <= 32'h1C003F00;
                                      char44_0[38] <= 32'h3C003F00;
                                      char44_0[39] <= 32'h7FFFFFFE;
                                      char44_0[40] <= 32'h7FFFFFFE;
                                      char44_0[41] <= 32'h00003F00;
                                      char44_0[42] <= 32'h00003F00;
                                      char44_0[43] <= 32'h00003F00;
                                      char44_0[44] <= 32'h00003F00;
                                      char44_0[45] <= 32'h00003F00;
                                      char44_0[46] <= 32'h00003F00;
                                      char44_0[47] <= 32'h00003F00;
                                      char44_0[48] <= 32'h00003F00;
                                      char44_0[49] <= 32'h00003F00;
                                      char44_0[50] <= 32'h00003F00;
                                      char44_0[51] <= 32'h00007F80;
                                      char44_0[52] <= 32'h000FFFFC;
                                      char44_0[53] <= 32'h000FFFFC;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//4
                                  4'd5: begin
                                      char44_0[  0] <= 32'h00000000;
                                      char44_0[  1] <= 32'h00000000;
                                      char44_0[  2] <= 32'h00000000;
                                      char44_0[  3] <= 32'h00000000;
                                      char44_0[  4] <= 32'h00000000;
                                      char44_0[  5] <= 32'h00000000;
                                      char44_0[  6] <= 32'h00000000;
                                      char44_0[  7] <= 32'h00000000;
                                      char44_0[  8] <= 32'h00000000;
                                      char44_0[  9] <= 32'h00000000;
                                      char44_0[10] <= 32'h00000000;
                                      char44_0[11] <= 32'h03FFFFF0;
                                      char44_0[12] <= 32'h03FFFFF0;
                                      char44_0[13] <= 32'h03FFFFF0;
                                      char44_0[14] <= 32'h03FFFFE0;
                                      char44_0[15] <= 32'h03800000;
                                      char44_0[16] <= 32'h03800000;
                                      char44_0[17] <= 32'h03800000;
                                      char44_0[18] <= 32'h03800000;
                                      char44_0[19] <= 32'h03800000;
                                      char44_0[20] <= 32'h07800000;
                                      char44_0[21] <= 32'h07800000;
                                      char44_0[22] <= 32'h07800000;
                                      char44_0[23] <= 32'h07800000;
                                      char44_0[24] <= 32'h07800000;
                                      char44_0[25] <= 32'h07800000;
                                      char44_0[26] <= 32'h078FF800;
                                      char44_0[27] <= 32'h073FFE00;
                                      char44_0[28] <= 32'h077FFF80;
                                      char44_0[29] <= 32'h07FC3F80;
                                      char44_0[30] <= 32'h07E00FC0;
                                      char44_0[31] <= 32'h07C007E0;
                                      char44_0[32] <= 32'h078007E0;
                                      char44_0[33] <= 32'h078003F0;
                                      char44_0[34] <= 32'h000003F0;
                                      char44_0[35] <= 32'h000001F0;
                                      char44_0[36] <= 32'h000001F8;
                                      char44_0[37] <= 32'h000001F8;
                                      char44_0[38] <= 32'h000001F8;
                                      char44_0[39] <= 32'h000001F8;
                                      char44_0[40] <= 32'h000001F8;
                                      char44_0[41] <= 32'h078001F8;
                                      char44_0[42] <= 32'h0FC001F8;
                                      char44_0[43] <= 32'h1FC001F0;
                                      char44_0[44] <= 32'h1FC001F0;
                                      char44_0[45] <= 32'h1FC003F0;
                                      char44_0[46] <= 32'h1F8003F0;
                                      char44_0[47] <= 32'h1F8003E0;
                                      char44_0[48] <= 32'h0F8007E0;
                                      char44_0[49] <= 32'h078007C0;
                                      char44_0[50] <= 32'h07C01F80;
                                      char44_0[51] <= 32'h03F83F00;
                                      char44_0[52] <= 32'h00FFFE00;
                                      char44_0[53] <= 32'h003FF800;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//5
                                  4'd6: begin
                                      char44_0[0] <= 32'h00000000;
                                      char44_0[1] <= 32'h00000000;
                                      char44_0[2] <= 32'h00000000;
                                      char44_0[3] <= 32'h00000000;
                                      char44_0[4] <= 32'h00000000;
                                      char44_0[5] <= 32'h00000000;
                                      char44_0[6] <= 32'h00000000;
                                      char44_0[7] <= 32'h00000000;
                                      char44_0[8] <= 32'h00000000;
                                      char44_0[9] <= 32'h00000000;
                                      char44_0[10] <= 32'h0007FE00;
                                      char44_0[11] <= 32'h001FFF80;
                                      char44_0[12] <= 32'h003F0FC0;
                                      char44_0[13] <= 32'h007C07C0;
                                      char44_0[14] <= 32'h00F807E0;
                                      char44_0[15] <= 32'h01F007E0;
                                      char44_0[16] <= 32'h03E007E0;
                                      char44_0[17] <= 32'h03C007E0;
                                      char44_0[18] <= 32'h07C003C0;
                                      char44_0[19] <= 32'h07C00000;
                                      char44_0[20] <= 32'h0FC00000;
                                      char44_0[21] <= 32'h0F800000;
                                      char44_0[22] <= 32'h0F800000;
                                      char44_0[23] <= 32'h1F800000;
                                      char44_0[24] <= 32'h1F800000;
                                      char44_0[25] <= 32'h1F800000;
                                      char44_0[26] <= 32'h1F87FE00;
                                      char44_0[27] <= 32'h1F9FFF80;
                                      char44_0[28] <= 32'h1FBFFFC0;
                                      char44_0[29] <= 32'h3FFE1FC0;
                                      char44_0[30] <= 32'h3FF807E0;
                                      char44_0[31] <= 32'h3FE003F0;
                                      char44_0[32] <= 32'h3FE003F0;
                                      char44_0[33] <= 32'h3FC001F8;
                                      char44_0[34] <= 32'h3F8001F8;
                                      char44_0[35] <= 32'h3F8001F8;
                                      char44_0[36] <= 32'h3F8000F8;
                                      char44_0[37] <= 32'h3F8000F8;
                                      char44_0[38] <= 32'h3F8000F8;
                                      char44_0[39] <= 32'h1F8000F8;
                                      char44_0[40] <= 32'h1F8000F8;
                                      char44_0[41] <= 32'h1F8000F8;
                                      char44_0[42] <= 32'h1F8000F8;
                                      char44_0[43] <= 32'h1F8000F8;
                                      char44_0[44] <= 32'h0FC001F8;
                                      char44_0[45] <= 32'h0FC001F8;
                                      char44_0[46] <= 32'h0FC001F0;
                                      char44_0[47] <= 32'h07E001F0;
                                      char44_0[48] <= 32'h03E003E0;
                                      char44_0[49] <= 32'h03F003E0;
                                      char44_0[50] <= 32'h01F807C0;
                                      char44_0[51] <= 32'h00FE1F80;
                                      char44_0[52] <= 32'h007FFE00;
                                      char44_0[53] <= 32'h001FF800;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//6
                                  4'd7: begin
                                      char44_0[0] <= 32'h00000000;
                                      char44_0[1] <= 32'h00000000;
                                      char44_0[2] <= 32'h00000000;
                                      char44_0[3] <= 32'h00000000;
                                      char44_0[4] <= 32'h00000000;
                                      char44_0[5] <= 32'h00000000;
                                      char44_0[6] <= 32'h00000000;
                                      char44_0[7] <= 32'h00000000;
                                      char44_0[8] <= 32'h00000000;
                                      char44_0[9] <= 32'h00000000;
                                      char44_0[10] <= 32'h00000000;
                                      char44_0[11] <= 32'h07FFFFF8;
                                      char44_0[12] <= 32'h07FFFFF8;
                                      char44_0[13] <= 32'h07FFFFF8;
                                      char44_0[14] <= 32'h0FFFFFF0;
                                      char44_0[15] <= 32'h0FC000E0;
                                      char44_0[16] <= 32'h0F8001E0;
                                      char44_0[17] <= 32'h0F0001C0;
                                      char44_0[18] <= 32'h0E0003C0;
                                      char44_0[19] <= 32'h0E000780;
                                      char44_0[20] <= 32'h1E000780;
                                      char44_0[21] <= 32'h1C000F00;
                                      char44_0[22] <= 32'h00000F00;
                                      char44_0[23] <= 32'h00001E00;
                                      char44_0[24] <= 32'h00001E00;
                                      char44_0[25] <= 32'h00003C00;
                                      char44_0[26] <= 32'h00003C00;
                                      char44_0[27] <= 32'h00007800;
                                      char44_0[28] <= 32'h00007800;
                                      char44_0[29] <= 32'h0000F800;
                                      char44_0[30] <= 32'h0000F000;
                                      char44_0[31] <= 32'h0001F000;
                                      char44_0[32] <= 32'h0001E000;
                                      char44_0[33] <= 32'h0003E000;
                                      char44_0[34] <= 32'h0003E000;
                                      char44_0[35] <= 32'h0003E000;
                                      char44_0[36] <= 32'h0007C000;
                                      char44_0[37] <= 32'h0007C000;
                                      char44_0[38] <= 32'h0007C000;
                                      char44_0[39] <= 32'h000FC000;
                                      char44_0[40] <= 32'h000FC000;
                                      char44_0[41] <= 32'h000FC000;
                                      char44_0[42] <= 32'h000FC000;
                                      char44_0[43] <= 32'h001FC000;
                                      char44_0[44] <= 32'h001FC000;
                                      char44_0[45] <= 32'h001FC000;
                                      char44_0[46] <= 32'h001FC000;
                                      char44_0[47] <= 32'h001FC000;
                                      char44_0[48] <= 32'h001FC000;
                                      char44_0[49] <= 32'h001FC000;
                                      char44_0[50] <= 32'h001FC000;
                                      char44_0[51] <= 32'h001FC000;
                                      char44_0[52] <= 32'h001FC000;
                                      char44_0[53] <= 32'h000F8000;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//7
                                  4'd8: begin
                                      char44_0[0] <= 32'h00000000;
                                      char44_0[1] <= 32'h00000000;
                                      char44_0[2] <= 32'h00000000;
                                      char44_0[3] <= 32'h00000000;
                                      char44_0[4] <= 32'h00000000;
                                      char44_0[5] <= 32'h00000000;
                                      char44_0[6] <= 32'h00000000;
                                      char44_0[7] <= 32'h00000000;
                                      char44_0[8] <= 32'h00000000;
                                      char44_0[9] <= 32'h00000000;
                                      char44_0[10] <= 32'h003FF800;
                                      char44_0[11] <= 32'h00FFFE00;
                                      char44_0[12] <= 32'h01F81F80;
                                      char44_0[13] <= 32'h03E00FC0;
                                      char44_0[14] <= 32'h07C003E0;
                                      char44_0[15] <= 32'h0F8003E0;
                                      char44_0[16] <= 32'h0F8001F0;
                                      char44_0[17] <= 32'h1F0001F0;
                                      char44_0[18] <= 32'h1F0001F0;
                                      char44_0[19] <= 32'h1F0001F0;
                                      char44_0[20] <= 32'h1F0001F0;
                                      char44_0[21] <= 32'h1F0001F0;
                                      char44_0[22] <= 32'h1F8001F0;
                                      char44_0[23] <= 32'h1FC001F0;
                                      char44_0[24] <= 32'h0FC001F0;
                                      char44_0[25] <= 32'h0FF003E0;
                                      char44_0[26] <= 32'h07F803C0;
                                      char44_0[27] <= 32'h03FE0F80;
                                      char44_0[28] <= 32'h01FF9F00;
                                      char44_0[29] <= 32'h00FFFE00;
                                      char44_0[30] <= 32'h003FF800;
                                      char44_0[31] <= 32'h007FFC00;
                                      char44_0[32] <= 32'h01F7FF00;
                                      char44_0[33] <= 32'h03E1FF80;
                                      char44_0[34] <= 32'h07C07FC0;
                                      char44_0[35] <= 32'h0F801FE0;
                                      char44_0[36] <= 32'h0F800FE0;
                                      char44_0[37] <= 32'h1F0007F0;
                                      char44_0[38] <= 32'h1F0003F0;
                                      char44_0[39] <= 32'h3E0001F8;
                                      char44_0[40] <= 32'h3E0001F8;
                                      char44_0[41] <= 32'h3E0001F8;
                                      char44_0[42] <= 32'h3E0000F8;
                                      char44_0[43] <= 32'h3E0000F8;
                                      char44_0[44] <= 32'h3E0000F8;
                                      char44_0[45] <= 32'h3E0000F8;
                                      char44_0[46] <= 32'h1F0001F0;
                                      char44_0[47] <= 32'h1F0001F0;
                                      char44_0[48] <= 32'h0F8003E0;
                                      char44_0[49] <= 32'h0FC003E0;
                                      char44_0[50] <= 32'h07E007C0;
                                      char44_0[51] <= 32'h01F83F80;
                                      char44_0[52] <= 32'h00FFFE00;
                                      char44_0[53] <= 32'h003FF800;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//8
                                  4'd9: begin
                                      char44_0[0] <= 32'h00000000;
                                      char44_0[1] <= 32'h00000000;
                                      char44_0[2] <= 32'h00000000;
                                      char44_0[3] <= 32'h00000000;
                                      char44_0[4] <= 32'h00000000;
                                      char44_0[5] <= 32'h00000000;
                                      char44_0[6] <= 32'h00000000;
                                      char44_0[7] <= 32'h00000000;
                                      char44_0[8] <= 32'h00000000;
                                      char44_0[9] <= 32'h00000000;
                                      char44_0[10] <= 32'h003FF000;
                                      char44_0[11] <= 32'h00FFFC00;
                                      char44_0[12] <= 32'h01F83F00;
                                      char44_0[13] <= 32'h03E01F80;
                                      char44_0[14] <= 32'h07C00F80;
                                      char44_0[15] <= 32'h0FC007C0;
                                      char44_0[16] <= 32'h0F8003E0;
                                      char44_0[17] <= 32'h1F8003E0;
                                      char44_0[18] <= 32'h1F0003F0;
                                      char44_0[19] <= 32'h1F0003F0;
                                      char44_0[20] <= 32'h3F0001F0;
                                      char44_0[21] <= 32'h3F0001F0;
                                      char44_0[22] <= 32'h3F0001F8;
                                      char44_0[23] <= 32'h3F0001F8;
                                      char44_0[24] <= 32'h3F0001F8;
                                      char44_0[25] <= 32'h3F0001F8;
                                      char44_0[26] <= 32'h3F0001F8;
                                      char44_0[27] <= 32'h3F0001F8;
                                      char44_0[28] <= 32'h3F0003F8;
                                      char44_0[29] <= 32'h1F8003F8;
                                      char44_0[30] <= 32'h1F8007F8;
                                      char44_0[31] <= 32'h1F800FF8;
                                      char44_0[32] <= 32'h0FC01FF8;
                                      char44_0[33] <= 32'h0FE03FF8;
                                      char44_0[34] <= 32'h07F8FDF8;
                                      char44_0[35] <= 32'h03FFF9F8;
                                      char44_0[36] <= 32'h01FFF1F8;
                                      char44_0[37] <= 32'h003F83F8;
                                      char44_0[38] <= 32'h000003F0;
                                      char44_0[39] <= 32'h000003F0;
                                      char44_0[40] <= 32'h000003F0;
                                      char44_0[41] <= 32'h000003F0;
                                      char44_0[42] <= 32'h000007E0;
                                      char44_0[43] <= 32'h000007E0;
                                      char44_0[44] <= 32'h000007C0;
                                      char44_0[45] <= 32'h03C007C0;
                                      char44_0[46] <= 32'h07C00F80;
                                      char44_0[47] <= 32'h0FE00F80;
                                      char44_0[48] <= 32'h0FE01F00;
                                      char44_0[49] <= 32'h0FE03E00;
                                      char44_0[50] <= 32'h07E07E00;
                                      char44_0[51] <= 32'h07F1F800;
                                      char44_0[52] <= 32'h03FFF000;
                                      char44_0[53] <= 32'h00FFC000;
                                      char44_0[54] <= 32'h00000000;
                                      char44_0[55] <= 32'h00000000;
                                      char44_0[56] <= 32'h00000000;
                                      char44_0[57] <= 32'h00000000;
                                      char44_0[58] <= 32'h00000000;
                                      char44_0[59] <= 32'h00000000;
                                      char44_0[60] <= 32'h00000000;
                                      char44_0[61] <= 32'h00000000;
                                      char44_0[62] <= 32'h00000000;
                                      char44_0[63] <= 32'h00000000;
                                  end//9
                                  default: begin
                                      char44_0[0] <= char44_0[0];
                                      char44_0[1] <= char44_0[1];
                                      char44_0[2] <= char44_0[2];
                                      char44_0[3] <= char44_0[3];
                                      char44_0[4] <= char44_0[4];
                                      char44_0[5] <= char44_0[5];
                                      char44_0[6] <= char44_0[6];
                                      char44_0[7] <= char44_0[7];
                                      char44_0[8] <= char44_0[8];
                                      char44_0[9] <= char44_0[9];
                                      char44_0[10] <= char44_0[10];
                                      char44_0[11] <= char44_0[11];
                                      char44_0[12] <= char44_0[12];
                                      char44_0[13] <= char44_0[13];
                                      char44_0[14] <= char44_0[14];
                                      char44_0[15] <= char44_0[15];
                                      char44_0[16] <= char44_0[16];
                                      char44_0[17] <= char44_0[17];
                                      char44_0[18] <= char44_0[18];
                                      char44_0[19] <= char44_0[19];
                                      char44_0[20] <= char44_0[20];
                                      char44_0[21] <= char44_0[21];
                                      char44_0[22] <= char44_0[22];
                                      char44_0[23] <= char44_0[23];
                                      char44_0[24] <= char44_0[24];
                                      char44_0[25] <= char44_0[25];
                                      char44_0[26] <= char44_0[26];
                                      char44_0[27] <= char44_0[27];
                                      char44_0[28] <= char44_0[28];
                                      char44_0[29] <= char44_0[29];
                                      char44_0[30] <= char44_0[30];
                                      char44_0[31] <= char44_0[31];
                                      char44_0[32] <= char44_0[32];
                                      char44_0[33] <= char44_0[33];
                                      char44_0[34] <= char44_0[34];
                                      char44_0[35] <= char44_0[35];
                                      char44_0[36] <= char44_0[36];
                                      char44_0[37] <= char44_0[37];
                                      char44_0[38] <= char44_0[38];
                                      char44_0[39] <= char44_0[39];
                                      char44_0[40] <= char44_0[40];
                                      char44_0[41] <= char44_0[41];
                                      char44_0[42] <= char44_0[42];
                                      char44_0[43] <= char44_0[43];
                                      char44_0[44] <= char44_0[44];
                                      char44_0[45] <= char44_0[45];
                                      char44_0[46] <= char44_0[46];
                                      char44_0[47] <= char44_0[47];
                                      char44_0[48] <= char44_0[48];
                                      char44_0[49] <= char44_0[49];
                                      char44_0[50] <= char44_0[50];
                                      char44_0[51] <= char44_0[51];
                                      char44_0[52] <= char44_0[52];
                                      char44_0[53] <= char44_0[53];
                                      char44_0[54] <= char44_0[54];
                                      char44_0[55] <= char44_0[55];
                                      char44_0[56] <= char44_0[56];
                                      char44_0[57] <= char44_0[57];
                                      char44_0[58] <= char44_0[58];
                                      char44_0[59] <= char44_0[59];
                                      char44_0[60] <= char44_0[60];
                                      char44_0[61] <= char44_0[61];
                                      char44_0[62] <= char44_0[62];
                                      char44_0[63] <= char44_0[63];
                                  end
                              endcase
                          
                              case((a2 - w1*(a2/w1))/k1)
                                      4'd0: begin
                                          char44_1[  0] <= 32'h00000000;
                                          char44_1[  1] <= 32'h00000000;
                                          char44_1[  2] <= 32'h00000000;
                                          char44_1[  3] <= 32'h00000000;
                                          char44_1[  4] <= 32'h00000000;
                                          char44_1[  5] <= 32'h00000000;
                                          char44_1[  6] <= 32'h00000000;
                                          char44_1[  7] <= 32'h00000000;
                                          char44_1[  8] <= 32'h00000000;
                                          char44_1[  9] <= 32'h00000000;
                                          char44_1[10] <= 32'h000FF000;
                                          char44_1[11] <= 32'h003FFC00;
                                          char44_1[12] <= 32'h007E7E00;
                                          char44_1[13] <= 32'h00F81F00;
                                          char44_1[14] <= 32'h01F00F80;
                                          char44_1[15] <= 32'h03F00FC0;
                                          char44_1[16] <= 32'h03E007C0;
                                          char44_1[17] <= 32'h07E007E0;
                                          char44_1[18] <= 32'h07C003E0;
                                          char44_1[19] <= 32'h0FC003F0;
                                          char44_1[20] <= 32'h0FC003F0;
                                          char44_1[21] <= 32'h0FC003F0;
                                          char44_1[22] <= 32'h1F8001F8;
                                          char44_1[23] <= 32'h1F8001F8;
                                          char44_1[24] <= 32'h1F8001F8;
                                          char44_1[25] <= 32'h1F8001F8;
                                          char44_1[26] <= 32'h1F8001F8;
                                          char44_1[27] <= 32'h3F8001F8;
                                          char44_1[28] <= 32'h3F8001F8;
                                          char44_1[29] <= 32'h3F8001F8;
                                          char44_1[30] <= 32'h3F8001F8;
                                          char44_1[31] <= 32'h3F8001F8;
                                          char44_1[32] <= 32'h3F8001F8;
                                          char44_1[33] <= 32'h3F8001F8;
                                          char44_1[34] <= 32'h3F8001F8;
                                          char44_1[35] <= 32'h3F8001F8;
                                          char44_1[36] <= 32'h3F8001F8;
                                          char44_1[37] <= 32'h1F8001F8;
                                          char44_1[38] <= 32'h1F8001F8;
                                          char44_1[39] <= 32'h1F8001F8;
                                          char44_1[40] <= 32'h1F8001F8;
                                          char44_1[41] <= 32'h1F8001F0;
                                          char44_1[42] <= 32'h0F8003F0;
                                          char44_1[43] <= 32'h0FC003F0;
                                          char44_1[44] <= 32'h0FC003F0;
                                          char44_1[45] <= 32'h07C003E0;
                                          char44_1[46] <= 32'h07E007E0;
                                          char44_1[47] <= 32'h03E007C0;
                                          char44_1[48] <= 32'h03F00FC0;
                                          char44_1[49] <= 32'h01F00F80;
                                          char44_1[50] <= 32'h00F81F00;
                                          char44_1[51] <= 32'h007E7E00;
                                          char44_1[52] <= 32'h003FFC00;
                                          char44_1[53] <= 32'h000FF000;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//0
                                      4'd1: begin
                                          char44_1[  0] <= 32'h00000000;
                                          char44_1[  1] <= 32'h00000000;
                                          char44_1[  2] <= 32'h00000000;
                                          char44_1[  3] <= 32'h00000000;
                                          char44_1[  4] <= 32'h00000000;
                                          char44_1[  5] <= 32'h00000000;
                                          char44_1[  6] <= 32'h00000000;
                                          char44_1[  7] <= 32'h00000000;
                                          char44_1[  8] <= 32'h00000000;
                                          char44_1[  9] <= 32'h00000000;
                                          char44_1[10] <= 32'h0000E000;
                                          char44_1[11] <= 32'h0001E000;
                                          char44_1[12] <= 32'h0003E000;
                                          char44_1[13] <= 32'h001FE000;
                                          char44_1[14] <= 32'h03FFE000;
                                          char44_1[15] <= 32'h03FFE000;
                                          char44_1[16] <= 32'h0007E000;
                                          char44_1[17] <= 32'h0007E000;
                                          char44_1[18] <= 32'h0007E000;
                                          char44_1[19] <= 32'h0007E000;
                                          char44_1[20] <= 32'h0007E000;
                                          char44_1[21] <= 32'h0007E000;
                                          char44_1[22] <= 32'h0007E000;
                                          char44_1[23] <= 32'h0007E000;
                                          char44_1[24] <= 32'h0007E000;
                                          char44_1[25] <= 32'h0007E000;
                                          char44_1[26] <= 32'h0007E000;
                                          char44_1[27] <= 32'h0007E000;
                                          char44_1[28] <= 32'h0007E000;
                                          char44_1[29] <= 32'h0007E000;
                                          char44_1[30] <= 32'h0007E000;
                                          char44_1[31] <= 32'h0007E000;
                                          char44_1[32] <= 32'h0007E000;
                                          char44_1[33] <= 32'h0007E000;
                                          char44_1[34] <= 32'h0007E000;
                                          char44_1[35] <= 32'h0007E000;
                                          char44_1[36] <= 32'h0007E000;
                                          char44_1[37] <= 32'h0007E000;
                                          char44_1[38] <= 32'h0007E000;
                                          char44_1[39] <= 32'h0007E000;
                                          char44_1[40] <= 32'h0007E000;
                                          char44_1[41] <= 32'h0007E000;
                                          char44_1[42] <= 32'h0007E000;
                                          char44_1[43] <= 32'h0007E000;
                                          char44_1[44] <= 32'h0007E000;
                                          char44_1[45] <= 32'h0007E000;
                                          char44_1[46] <= 32'h0007E000;
                                          char44_1[47] <= 32'h0007E000;
                                          char44_1[48] <= 32'h0007E000;
                                          char44_1[49] <= 32'h0007E000;
                                          char44_1[50] <= 32'h0007E000;
                                          char44_1[51] <= 32'h000FF800;
                                          char44_1[52] <= 32'h03FFFFC0;
                                          char44_1[53] <= 32'h03FFFFC0;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//1
                                      4'd2: begin
                                          char44_1[  0] <= 32'h00000000;
                                          char44_1[  1] <= 32'h00000000;
                                          char44_1[  2] <= 32'h00000000;
                                          char44_1[  3] <= 32'h00000000;
                                          char44_1[  4] <= 32'h00000000;
                                          char44_1[  5] <= 32'h00000000;
                                          char44_1[  6] <= 32'h00000000;
                                          char44_1[  7] <= 32'h00000000;
                                          char44_1[  8] <= 32'h00000000;
                                          char44_1[  9] <= 32'h00000000;
                                          char44_1[10] <= 32'h001FFC00;
                                          char44_1[11] <= 32'h007FFF00;
                                          char44_1[12] <= 32'h01F83F80;
                                          char44_1[13] <= 32'h03E00FC0;
                                          char44_1[14] <= 32'h07C007E0;
                                          char44_1[15] <= 32'h078007E0;
                                          char44_1[16] <= 32'h0F8003F0;
                                          char44_1[17] <= 32'h0F8003F0;
                                          char44_1[18] <= 32'h1F8003F0;
                                          char44_1[19] <= 32'h1F8003F0;
                                          char44_1[20] <= 32'h1FC003F0;
                                          char44_1[21] <= 32'h1FC003F0;
                                          char44_1[22] <= 32'h1FC003F0;
                                          char44_1[23] <= 32'h0FC003F0;
                                          char44_1[24] <= 32'h07C003F0;
                                          char44_1[25] <= 32'h000003E0;
                                          char44_1[26] <= 32'h000007E0;
                                          char44_1[27] <= 32'h000007E0;
                                          char44_1[28] <= 32'h00000FC0;
                                          char44_1[29] <= 32'h00000F80;
                                          char44_1[30] <= 32'h00001F80;
                                          char44_1[31] <= 32'h00003F00;
                                          char44_1[32] <= 32'h00003E00;
                                          char44_1[33] <= 32'h00007C00;
                                          char44_1[34] <= 32'h0000F800;
                                          char44_1[35] <= 32'h0001F000;
                                          char44_1[36] <= 32'h0003E000;
                                          char44_1[37] <= 32'h0007C000;
                                          char44_1[38] <= 32'h000F8000;
                                          char44_1[39] <= 32'h001F0000;
                                          char44_1[40] <= 32'h003E0000;
                                          char44_1[41] <= 32'h007C0000;
                                          char44_1[42] <= 32'h00F80000;
                                          char44_1[43] <= 32'h01F00038;
                                          char44_1[44] <= 32'h01E00038;
                                          char44_1[45] <= 32'h03C00070;
                                          char44_1[46] <= 32'h07800070;
                                          char44_1[47] <= 32'h0F8000F0;
                                          char44_1[48] <= 32'h0F0000F0;
                                          char44_1[49] <= 32'h1E0003F0;
                                          char44_1[50] <= 32'h3FFFFFF0;
                                          char44_1[51] <= 32'h3FFFFFF0;
                                          char44_1[52] <= 32'h3FFFFFE0;
                                          char44_1[53] <= 32'h3FFFFFE0;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//2
                                      4'd3: begin
                                          char44_1[  0] <= 32'h00000000;
                                          char44_1[  1] <= 32'h00000000;
                                          char44_1[  2] <= 32'h00000000;
                                          char44_1[  3] <= 32'h00000000;
                                          char44_1[  4] <= 32'h00000000;
                                          char44_1[  5] <= 32'h00000000;
                                          char44_1[  6] <= 32'h00000000;
                                          char44_1[  7] <= 32'h00000000;
                                          char44_1[  8] <= 32'h00000000;
                                          char44_1[  9] <= 32'h00000000;
                                          char44_1[10] <= 32'h003FF000;
                                          char44_1[11] <= 32'h00FFFC00;
                                          char44_1[12] <= 32'h01F07E00;
                                          char44_1[13] <= 32'h03C03F00;
                                          char44_1[14] <= 32'h07801F80;
                                          char44_1[15] <= 32'h0F800FC0;
                                          char44_1[16] <= 32'h0F800FC0;
                                          char44_1[17] <= 32'h0F8007E0;
                                          char44_1[18] <= 32'h0FC007E0;
                                          char44_1[19] <= 32'h0FC007E0;
                                          char44_1[20] <= 32'h0FC007E0;
                                          char44_1[21] <= 32'h07C007E0;
                                          char44_1[22] <= 32'h000007E0;
                                          char44_1[23] <= 32'h000007E0;
                                          char44_1[24] <= 32'h000007C0;
                                          char44_1[25] <= 32'h00000FC0;
                                          char44_1[26] <= 32'h00000F80;
                                          char44_1[27] <= 32'h00001F00;
                                          char44_1[28] <= 32'h00007E00;
                                          char44_1[29] <= 32'h0003FC00;
                                          char44_1[30] <= 32'h001FF000;
                                          char44_1[31] <= 32'h001FFC00;
                                          char44_1[32] <= 32'h0000FF00;
                                          char44_1[33] <= 32'h00001F80;
                                          char44_1[34] <= 32'h00000FC0;
                                          char44_1[35] <= 32'h000007E0;
                                          char44_1[36] <= 32'h000003E0;
                                          char44_1[37] <= 32'h000003F0;
                                          char44_1[38] <= 32'h000003F0;
                                          char44_1[39] <= 32'h000001F0;
                                          char44_1[40] <= 32'h000001F8;
                                          char44_1[41] <= 32'h000001F8;
                                          char44_1[42] <= 32'h078001F8;
                                          char44_1[43] <= 32'h0FC001F8;
                                          char44_1[44] <= 32'h1FC001F8;
                                          char44_1[45] <= 32'h1FC003F0;
                                          char44_1[46] <= 32'h1FC003F0;
                                          char44_1[47] <= 32'h1FC003E0;
                                          char44_1[48] <= 32'h0F8007E0;
                                          char44_1[49] <= 32'h0F8007C0;
                                          char44_1[50] <= 32'h07C01F80;
                                          char44_1[51] <= 32'h03F07F00;
                                          char44_1[52] <= 32'h01FFFE00;
                                          char44_1[53] <= 32'h003FF000;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//3
                                      4'd4: begin
                                          char44_1[  0] <= 32'h00000000;
                                          char44_1[  1] <= 32'h00000000;
                                          char44_1[  2] <= 32'h00000000;
                                          char44_1[  3] <= 32'h00000000;
                                          char44_1[  4] <= 32'h00000000;
                                          char44_1[  5] <= 32'h00000000;
                                          char44_1[  6] <= 32'h00000000;
                                          char44_1[  7] <= 32'h00000000;
                                          char44_1[  8] <= 32'h00000000;
                                          char44_1[  9] <= 32'h00000000;
                                          char44_1[10] <= 32'h00001F00;
                                          char44_1[11] <= 32'h00001F00;
                                          char44_1[12] <= 32'h00003F00;
                                          char44_1[13] <= 32'h00003F00;
                                          char44_1[14] <= 32'h00007F00;
                                          char44_1[15] <= 32'h0000FF00;
                                          char44_1[16] <= 32'h0000FF00;
                                          char44_1[17] <= 32'h0001FF00;
                                          char44_1[18] <= 32'h0003FF00;
                                          char44_1[19] <= 32'h0003BF00;
                                          char44_1[20] <= 32'h0007BF00;
                                          char44_1[21] <= 32'h00073F00;
                                          char44_1[22] <= 32'h000F3F00;
                                          char44_1[23] <= 32'h001E3F00;
                                          char44_1[24] <= 32'h001C3F00;
                                          char44_1[25] <= 32'h003C3F00;
                                          char44_1[26] <= 32'h00783F00;
                                          char44_1[27] <= 32'h00783F00;
                                          char44_1[28] <= 32'h00F03F00;
                                          char44_1[29] <= 32'h00E03F00;
                                          char44_1[30] <= 32'h01E03F00;
                                          char44_1[31] <= 32'h03C03F00;
                                          char44_1[32] <= 32'h03803F00;
                                          char44_1[33] <= 32'h07803F00;
                                          char44_1[34] <= 32'h0F003F00;
                                          char44_1[35] <= 32'h0F003F00;
                                          char44_1[36] <= 32'h1E003F00;
                                          char44_1[37] <= 32'h1C003F00;
                                          char44_1[38] <= 32'h3C003F00;
                                          char44_1[39] <= 32'h7FFFFFFE;
                                          char44_1[40] <= 32'h7FFFFFFE;
                                          char44_1[41] <= 32'h00003F00;
                                          char44_1[42] <= 32'h00003F00;
                                          char44_1[43] <= 32'h00003F00;
                                          char44_1[44] <= 32'h00003F00;
                                          char44_1[45] <= 32'h00003F00;
                                          char44_1[46] <= 32'h00003F00;
                                          char44_1[47] <= 32'h00003F00;
                                          char44_1[48] <= 32'h00003F00;
                                          char44_1[49] <= 32'h00003F00;
                                          char44_1[50] <= 32'h00003F00;
                                          char44_1[51] <= 32'h00007F80;
                                          char44_1[52] <= 32'h000FFFFC;
                                          char44_1[53] <= 32'h000FFFFC;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//4
                                      4'd5: begin
                                          char44_1[  0] <= 32'h00000000;
                                          char44_1[  1] <= 32'h00000000;
                                          char44_1[  2] <= 32'h00000000;
                                          char44_1[  3] <= 32'h00000000;
                                          char44_1[  4] <= 32'h00000000;
                                          char44_1[  5] <= 32'h00000000;
                                          char44_1[  6] <= 32'h00000000;
                                          char44_1[  7] <= 32'h00000000;
                                          char44_1[  8] <= 32'h00000000;
                                          char44_1[  9] <= 32'h00000000;
                                          char44_1[10] <= 32'h00000000;
                                          char44_1[11] <= 32'h03FFFFF0;
                                          char44_1[12] <= 32'h03FFFFF0;
                                          char44_1[13] <= 32'h03FFFFF0;
                                          char44_1[14] <= 32'h03FFFFE0;
                                          char44_1[15] <= 32'h03800000;
                                          char44_1[16] <= 32'h03800000;
                                          char44_1[17] <= 32'h03800000;
                                          char44_1[18] <= 32'h03800000;
                                          char44_1[19] <= 32'h03800000;
                                          char44_1[20] <= 32'h07800000;
                                          char44_1[21] <= 32'h07800000;
                                          char44_1[22] <= 32'h07800000;
                                          char44_1[23] <= 32'h07800000;
                                          char44_1[24] <= 32'h07800000;
                                          char44_1[25] <= 32'h07800000;
                                          char44_1[26] <= 32'h078FF800;
                                          char44_1[27] <= 32'h073FFE00;
                                          char44_1[28] <= 32'h077FFF80;
                                          char44_1[29] <= 32'h07FC3F80;
                                          char44_1[30] <= 32'h07E00FC0;
                                          char44_1[31] <= 32'h07C007E0;
                                          char44_1[32] <= 32'h078007E0;
                                          char44_1[33] <= 32'h078003F0;
                                          char44_1[34] <= 32'h000003F0;
                                          char44_1[35] <= 32'h000001F0;
                                          char44_1[36] <= 32'h000001F8;
                                          char44_1[37] <= 32'h000001F8;
                                          char44_1[38] <= 32'h000001F8;
                                          char44_1[39] <= 32'h000001F8;
                                          char44_1[40] <= 32'h000001F8;
                                          char44_1[41] <= 32'h078001F8;
                                          char44_1[42] <= 32'h0FC001F8;
                                          char44_1[43] <= 32'h1FC001F0;
                                          char44_1[44] <= 32'h1FC001F0;
                                          char44_1[45] <= 32'h1FC003F0;
                                          char44_1[46] <= 32'h1F8003F0;
                                          char44_1[47] <= 32'h1F8003E0;
                                          char44_1[48] <= 32'h0F8007E0;
                                          char44_1[49] <= 32'h078007C0;
                                          char44_1[50] <= 32'h07C01F80;
                                          char44_1[51] <= 32'h03F83F00;
                                          char44_1[52] <= 32'h00FFFE00;
                                          char44_1[53] <= 32'h003FF800;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//5
                                      4'd6: begin
                                          char44_1[0] <= 32'h00000000;
                                          char44_1[1] <= 32'h00000000;
                                          char44_1[2] <= 32'h00000000;
                                          char44_1[3] <= 32'h00000000;
                                          char44_1[4] <= 32'h00000000;
                                          char44_1[5] <= 32'h00000000;
                                          char44_1[6] <= 32'h00000000;
                                          char44_1[7] <= 32'h00000000;
                                          char44_1[8] <= 32'h00000000;
                                          char44_1[9] <= 32'h00000000;
                                          char44_1[10] <= 32'h0007FE00;
                                          char44_1[11] <= 32'h001FFF80;
                                          char44_1[12] <= 32'h003F0FC0;
                                          char44_1[13] <= 32'h007C07C0;
                                          char44_1[14] <= 32'h00F807E0;
                                          char44_1[15] <= 32'h01F007E0;
                                          char44_1[16] <= 32'h03E007E0;
                                          char44_1[17] <= 32'h03C007E0;
                                          char44_1[18] <= 32'h07C003C0;
                                          char44_1[19] <= 32'h07C00000;
                                          char44_1[20] <= 32'h0FC00000;
                                          char44_1[21] <= 32'h0F800000;
                                          char44_1[22] <= 32'h0F800000;
                                          char44_1[23] <= 32'h1F800000;
                                          char44_1[24] <= 32'h1F800000;
                                          char44_1[25] <= 32'h1F800000;
                                          char44_1[26] <= 32'h1F87FE00;
                                          char44_1[27] <= 32'h1F9FFF80;
                                          char44_1[28] <= 32'h1FBFFFC0;
                                          char44_1[29] <= 32'h3FFE1FC0;
                                          char44_1[30] <= 32'h3FF807E0;
                                          char44_1[31] <= 32'h3FE003F0;
                                          char44_1[32] <= 32'h3FE003F0;
                                          char44_1[33] <= 32'h3FC001F8;
                                          char44_1[34] <= 32'h3F8001F8;
                                          char44_1[35] <= 32'h3F8001F8;
                                          char44_1[36] <= 32'h3F8000F8;
                                          char44_1[37] <= 32'h3F8000F8;
                                          char44_1[38] <= 32'h3F8000F8;
                                          char44_1[39] <= 32'h1F8000F8;
                                          char44_1[40] <= 32'h1F8000F8;
                                          char44_1[41] <= 32'h1F8000F8;
                                          char44_1[42] <= 32'h1F8000F8;
                                          char44_1[43] <= 32'h1F8000F8;
                                          char44_1[44] <= 32'h0FC001F8;
                                          char44_1[45] <= 32'h0FC001F8;
                                          char44_1[46] <= 32'h0FC001F0;
                                          char44_1[47] <= 32'h07E001F0;
                                          char44_1[48] <= 32'h03E003E0;
                                          char44_1[49] <= 32'h03F003E0;
                                          char44_1[50] <= 32'h01F807C0;
                                          char44_1[51] <= 32'h00FE1F80;
                                          char44_1[52] <= 32'h007FFE00;
                                          char44_1[53] <= 32'h001FF800;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//6
                                      4'd7: begin
                                          char44_1[0] <= 32'h00000000;
                                          char44_1[1] <= 32'h00000000;
                                          char44_1[2] <= 32'h00000000;
                                          char44_1[3] <= 32'h00000000;
                                          char44_1[4] <= 32'h00000000;
                                          char44_1[5] <= 32'h00000000;
                                          char44_1[6] <= 32'h00000000;
                                          char44_1[7] <= 32'h00000000;
                                          char44_1[8] <= 32'h00000000;
                                          char44_1[9] <= 32'h00000000;
                                          char44_1[10] <= 32'h00000000;
                                          char44_1[11] <= 32'h07FFFFF8;
                                          char44_1[12] <= 32'h07FFFFF8;
                                          char44_1[13] <= 32'h07FFFFF8;
                                          char44_1[14] <= 32'h0FFFFFF0;
                                          char44_1[15] <= 32'h0FC000E0;
                                          char44_1[16] <= 32'h0F8001E0;
                                          char44_1[17] <= 32'h0F0001C0;
                                          char44_1[18] <= 32'h0E0003C0;
                                          char44_1[19] <= 32'h0E000780;
                                          char44_1[20] <= 32'h1E000780;
                                          char44_1[21] <= 32'h1C000F00;
                                          char44_1[22] <= 32'h00000F00;
                                          char44_1[23] <= 32'h00001E00;
                                          char44_1[24] <= 32'h00001E00;
                                          char44_1[25] <= 32'h00003C00;
                                          char44_1[26] <= 32'h00003C00;
                                          char44_1[27] <= 32'h00007800;
                                          char44_1[28] <= 32'h00007800;
                                          char44_1[29] <= 32'h0000F800;
                                          char44_1[30] <= 32'h0000F000;
                                          char44_1[31] <= 32'h0001F000;
                                          char44_1[32] <= 32'h0001E000;
                                          char44_1[33] <= 32'h0003E000;
                                          char44_1[34] <= 32'h0003E000;
                                          char44_1[35] <= 32'h0003E000;
                                          char44_1[36] <= 32'h0007C000;
                                          char44_1[37] <= 32'h0007C000;
                                          char44_1[38] <= 32'h0007C000;
                                          char44_1[39] <= 32'h000FC000;
                                          char44_1[40] <= 32'h000FC000;
                                          char44_1[41] <= 32'h000FC000;
                                          char44_1[42] <= 32'h000FC000;
                                          char44_1[43] <= 32'h001FC000;
                                          char44_1[44] <= 32'h001FC000;
                                          char44_1[45] <= 32'h001FC000;
                                          char44_1[46] <= 32'h001FC000;
                                          char44_1[47] <= 32'h001FC000;
                                          char44_1[48] <= 32'h001FC000;
                                          char44_1[49] <= 32'h001FC000;
                                          char44_1[50] <= 32'h001FC000;
                                          char44_1[51] <= 32'h001FC000;
                                          char44_1[52] <= 32'h001FC000;
                                          char44_1[53] <= 32'h000F8000;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//7
                                      4'd8: begin
                                          char44_1[0] <= 32'h00000000;
                                          char44_1[1] <= 32'h00000000;
                                          char44_1[2] <= 32'h00000000;
                                          char44_1[3] <= 32'h00000000;
                                          char44_1[4] <= 32'h00000000;
                                          char44_1[5] <= 32'h00000000;
                                          char44_1[6] <= 32'h00000000;
                                          char44_1[7] <= 32'h00000000;
                                          char44_1[8] <= 32'h00000000;
                                          char44_1[9] <= 32'h00000000;
                                          char44_1[10] <= 32'h003FF800;
                                          char44_1[11] <= 32'h00FFFE00;
                                          char44_1[12] <= 32'h01F81F80;
                                          char44_1[13] <= 32'h03E00FC0;
                                          char44_1[14] <= 32'h07C003E0;
                                          char44_1[15] <= 32'h0F8003E0;
                                          char44_1[16] <= 32'h0F8001F0;
                                          char44_1[17] <= 32'h1F0001F0;
                                          char44_1[18] <= 32'h1F0001F0;
                                          char44_1[19] <= 32'h1F0001F0;
                                          char44_1[20] <= 32'h1F0001F0;
                                          char44_1[21] <= 32'h1F0001F0;
                                          char44_1[22] <= 32'h1F8001F0;
                                          char44_1[23] <= 32'h1FC001F0;
                                          char44_1[24] <= 32'h0FC001F0;
                                          char44_1[25] <= 32'h0FF003E0;
                                          char44_1[26] <= 32'h07F803C0;
                                          char44_1[27] <= 32'h03FE0F80;
                                          char44_1[28] <= 32'h01FF9F00;
                                          char44_1[29] <= 32'h00FFFE00;
                                          char44_1[30] <= 32'h003FF800;
                                          char44_1[31] <= 32'h007FFC00;
                                          char44_1[32] <= 32'h01F7FF00;
                                          char44_1[33] <= 32'h03E1FF80;
                                          char44_1[34] <= 32'h07C07FC0;
                                          char44_1[35] <= 32'h0F801FE0;
                                          char44_1[36] <= 32'h0F800FE0;
                                          char44_1[37] <= 32'h1F0007F0;
                                          char44_1[38] <= 32'h1F0003F0;
                                          char44_1[39] <= 32'h3E0001F8;
                                          char44_1[40] <= 32'h3E0001F8;
                                          char44_1[41] <= 32'h3E0001F8;
                                          char44_1[42] <= 32'h3E0000F8;
                                          char44_1[43] <= 32'h3E0000F8;
                                          char44_1[44] <= 32'h3E0000F8;
                                          char44_1[45] <= 32'h3E0000F8;
                                          char44_1[46] <= 32'h1F0001F0;
                                          char44_1[47] <= 32'h1F0001F0;
                                          char44_1[48] <= 32'h0F8003E0;
                                          char44_1[49] <= 32'h0FC003E0;
                                          char44_1[50] <= 32'h07E007C0;
                                          char44_1[51] <= 32'h01F83F80;
                                          char44_1[52] <= 32'h00FFFE00;
                                          char44_1[53] <= 32'h003FF800;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//8
                                      4'd9: begin
                                          char44_1[0] <= 32'h00000000;
                                          char44_1[1] <= 32'h00000000;
                                          char44_1[2] <= 32'h00000000;
                                          char44_1[3] <= 32'h00000000;
                                          char44_1[4] <= 32'h00000000;
                                          char44_1[5] <= 32'h00000000;
                                          char44_1[6] <= 32'h00000000;
                                          char44_1[7] <= 32'h00000000;
                                          char44_1[8] <= 32'h00000000;
                                          char44_1[9] <= 32'h00000000;
                                          char44_1[10] <= 32'h003FF000;
                                          char44_1[11] <= 32'h00FFFC00;
                                          char44_1[12] <= 32'h01F83F00;
                                          char44_1[13] <= 32'h03E01F80;
                                          char44_1[14] <= 32'h07C00F80;
                                          char44_1[15] <= 32'h0FC007C0;
                                          char44_1[16] <= 32'h0F8003E0;
                                          char44_1[17] <= 32'h1F8003E0;
                                          char44_1[18] <= 32'h1F0003F0;
                                          char44_1[19] <= 32'h1F0003F0;
                                          char44_1[20] <= 32'h3F0001F0;
                                          char44_1[21] <= 32'h3F0001F0;
                                          char44_1[22] <= 32'h3F0001F8;
                                          char44_1[23] <= 32'h3F0001F8;
                                          char44_1[24] <= 32'h3F0001F8;
                                          char44_1[25] <= 32'h3F0001F8;
                                          char44_1[26] <= 32'h3F0001F8;
                                          char44_1[27] <= 32'h3F0001F8;
                                          char44_1[28] <= 32'h3F0003F8;
                                          char44_1[29] <= 32'h1F8003F8;
                                          char44_1[30] <= 32'h1F8007F8;
                                          char44_1[31] <= 32'h1F800FF8;
                                          char44_1[32] <= 32'h0FC01FF8;
                                          char44_1[33] <= 32'h0FE03FF8;
                                          char44_1[34] <= 32'h07F8FDF8;
                                          char44_1[35] <= 32'h03FFF9F8;
                                          char44_1[36] <= 32'h01FFF1F8;
                                          char44_1[37] <= 32'h003F83F8;
                                          char44_1[38] <= 32'h000003F0;
                                          char44_1[39] <= 32'h000003F0;
                                          char44_1[40] <= 32'h000003F0;
                                          char44_1[41] <= 32'h000003F0;
                                          char44_1[42] <= 32'h000007E0;
                                          char44_1[43] <= 32'h000007E0;
                                          char44_1[44] <= 32'h000007C0;
                                          char44_1[45] <= 32'h03C007C0;
                                          char44_1[46] <= 32'h07C00F80;
                                          char44_1[47] <= 32'h0FE00F80;
                                          char44_1[48] <= 32'h0FE01F00;
                                          char44_1[49] <= 32'h0FE03E00;
                                          char44_1[50] <= 32'h07E07E00;
                                          char44_1[51] <= 32'h07F1F800;
                                          char44_1[52] <= 32'h03FFF000;
                                          char44_1[53] <= 32'h00FFC000;
                                          char44_1[54] <= 32'h00000000;
                                          char44_1[55] <= 32'h00000000;
                                          char44_1[56] <= 32'h00000000;
                                          char44_1[57] <= 32'h00000000;
                                          char44_1[58] <= 32'h00000000;
                                          char44_1[59] <= 32'h00000000;
                                          char44_1[60] <= 32'h00000000;
                                          char44_1[61] <= 32'h00000000;
                                          char44_1[62] <= 32'h00000000;
                                          char44_1[63] <= 32'h00000000;
                                      end//9
                                      default: begin
                                          char44_1[0] <= char44_1[0];
                                          char44_1[1] <= char44_1[1];
                                          char44_1[2] <= char44_1[2];
                                          char44_1[3] <= char44_1[3];
                                          char44_1[4] <= char44_1[4];
                                          char44_1[5] <= char44_1[5];
                                          char44_1[6] <= char44_1[6];
                                          char44_1[7] <= char44_1[7];
                                          char44_1[8] <= char44_1[8];
                                          char44_1[9] <= char44_1[9];
                                          char44_1[10] <= char44_1[10];
                                          char44_1[11] <= char44_1[11];
                                          char44_1[12] <= char44_1[12];
                                          char44_1[13] <= char44_1[13];
                                          char44_1[14] <= char44_1[14];
                                          char44_1[15] <= char44_1[15];
                                          char44_1[16] <= char44_1[16];
                                          char44_1[17] <= char44_1[17];
                                          char44_1[18] <= char44_1[18];
                                          char44_1[19] <= char44_1[19];
                                          char44_1[20] <= char44_1[20];
                                          char44_1[21] <= char44_1[21];
                                          char44_1[22] <= char44_1[22];
                                          char44_1[23] <= char44_1[23];
                                          char44_1[24] <= char44_1[24];
                                          char44_1[25] <= char44_1[25];
                                          char44_1[26] <= char44_1[26];
                                          char44_1[27] <= char44_1[27];
                                          char44_1[28] <= char44_1[28];
                                          char44_1[29] <= char44_1[29];
                                          char44_1[30] <= char44_1[30];
                                          char44_1[31] <= char44_1[31];
                                          char44_1[32] <= char44_1[32];
                                          char44_1[33] <= char44_1[33];
                                          char44_1[34] <= char44_1[34];
                                          char44_1[35] <= char44_1[35];
                                          char44_1[36] <= char44_1[36];
                                          char44_1[37] <= char44_1[37];
                                          char44_1[38] <= char44_1[38];
                                          char44_1[39] <= char44_1[39];
                                          char44_1[40] <= char44_1[40];
                                          char44_1[41] <= char44_1[41];
                                          char44_1[42] <= char44_1[42];
                                          char44_1[43] <= char44_1[43];
                                          char44_1[44] <= char44_1[44];
                                          char44_1[45] <= char44_1[45];
                                          char44_1[46] <= char44_1[46];
                                          char44_1[47] <= char44_1[47];
                                          char44_1[48] <= char44_1[48];
                                          char44_1[49] <= char44_1[49];
                                          char44_1[50] <= char44_1[50];
                                          char44_1[51] <= char44_1[51];
                                          char44_1[52] <= char44_1[52];
                                          char44_1[53] <= char44_1[53];
                                          char44_1[54] <= char44_1[54];
                                          char44_1[55] <= char44_1[55];
                                          char44_1[56] <= char44_1[56];
                                          char44_1[57] <= char44_1[57];
                                          char44_1[58] <= char44_1[58];
                                          char44_1[59] <= char44_1[59];
                                          char44_1[60] <= char44_1[60];
                                          char44_1[61] <= char44_1[61];
                                          char44_1[62] <= char44_1[62];
                                          char44_1[63] <= char44_1[63];
                                      end
                                  endcase
                          
                              case((a2 - k1*(a2/k1))/h1)
                                          4'd0: begin
                                              char44_2[  0] <= 32'h00000000;
                                              char44_2[  1] <= 32'h00000000;
                                              char44_2[  2] <= 32'h00000000;
                                              char44_2[  3] <= 32'h00000000;
                                              char44_2[  4] <= 32'h00000000;
                                              char44_2[  5] <= 32'h00000000;
                                              char44_2[  6] <= 32'h00000000;
                                              char44_2[  7] <= 32'h00000000;
                                              char44_2[  8] <= 32'h00000000;
                                              char44_2[  9] <= 32'h00000000;
                                              char44_2[10] <= 32'h000FF000;
                                              char44_2[11] <= 32'h003FFC00;
                                              char44_2[12] <= 32'h007E7E00;
                                              char44_2[13] <= 32'h00F81F00;
                                              char44_2[14] <= 32'h01F00F80;
                                              char44_2[15] <= 32'h03F00FC0;
                                              char44_2[16] <= 32'h03E007C0;
                                              char44_2[17] <= 32'h07E007E0;
                                              char44_2[18] <= 32'h07C003E0;
                                              char44_2[19] <= 32'h0FC003F0;
                                              char44_2[20] <= 32'h0FC003F0;
                                              char44_2[21] <= 32'h0FC003F0;
                                              char44_2[22] <= 32'h1F8001F8;
                                              char44_2[23] <= 32'h1F8001F8;
                                              char44_2[24] <= 32'h1F8001F8;
                                              char44_2[25] <= 32'h1F8001F8;
                                              char44_2[26] <= 32'h1F8001F8;
                                              char44_2[27] <= 32'h3F8001F8;
                                              char44_2[28] <= 32'h3F8001F8;
                                              char44_2[29] <= 32'h3F8001F8;
                                              char44_2[30] <= 32'h3F8001F8;
                                              char44_2[31] <= 32'h3F8001F8;
                                              char44_2[32] <= 32'h3F8001F8;
                                              char44_2[33] <= 32'h3F8001F8;
                                              char44_2[34] <= 32'h3F8001F8;
                                              char44_2[35] <= 32'h3F8001F8;
                                              char44_2[36] <= 32'h3F8001F8;
                                              char44_2[37] <= 32'h1F8001F8;
                                              char44_2[38] <= 32'h1F8001F8;
                                              char44_2[39] <= 32'h1F8001F8;
                                              char44_2[40] <= 32'h1F8001F8;
                                              char44_2[41] <= 32'h1F8001F0;
                                              char44_2[42] <= 32'h0F8003F0;
                                              char44_2[43] <= 32'h0FC003F0;
                                              char44_2[44] <= 32'h0FC003F0;
                                              char44_2[45] <= 32'h07C003E0;
                                              char44_2[46] <= 32'h07E007E0;
                                              char44_2[47] <= 32'h03E007C0;
                                              char44_2[48] <= 32'h03F00FC0;
                                              char44_2[49] <= 32'h01F00F80;
                                              char44_2[50] <= 32'h00F81F00;
                                              char44_2[51] <= 32'h007E7E00;
                                              char44_2[52] <= 32'h003FFC00;
                                              char44_2[53] <= 32'h000FF000;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//0
                                          4'd1: begin
                                              char44_2[  0] <= 32'h00000000;
                                              char44_2[  1] <= 32'h00000000;
                                              char44_2[  2] <= 32'h00000000;
                                              char44_2[  3] <= 32'h00000000;
                                              char44_2[  4] <= 32'h00000000;
                                              char44_2[  5] <= 32'h00000000;
                                              char44_2[  6] <= 32'h00000000;
                                              char44_2[  7] <= 32'h00000000;
                                              char44_2[  8] <= 32'h00000000;
                                              char44_2[  9] <= 32'h00000000;
                                              char44_2[10] <= 32'h0000E000;
                                              char44_2[11] <= 32'h0001E000;
                                              char44_2[12] <= 32'h0003E000;
                                              char44_2[13] <= 32'h001FE000;
                                              char44_2[14] <= 32'h03FFE000;
                                              char44_2[15] <= 32'h03FFE000;
                                              char44_2[16] <= 32'h0007E000;
                                              char44_2[17] <= 32'h0007E000;
                                              char44_2[18] <= 32'h0007E000;
                                              char44_2[19] <= 32'h0007E000;
                                              char44_2[20] <= 32'h0007E000;
                                              char44_2[21] <= 32'h0007E000;
                                              char44_2[22] <= 32'h0007E000;
                                              char44_2[23] <= 32'h0007E000;
                                              char44_2[24] <= 32'h0007E000;
                                              char44_2[25] <= 32'h0007E000;
                                              char44_2[26] <= 32'h0007E000;
                                              char44_2[27] <= 32'h0007E000;
                                              char44_2[28] <= 32'h0007E000;
                                              char44_2[29] <= 32'h0007E000;
                                              char44_2[30] <= 32'h0007E000;
                                              char44_2[31] <= 32'h0007E000;
                                              char44_2[32] <= 32'h0007E000;
                                              char44_2[33] <= 32'h0007E000;
                                              char44_2[34] <= 32'h0007E000;
                                              char44_2[35] <= 32'h0007E000;
                                              char44_2[36] <= 32'h0007E000;
                                              char44_2[37] <= 32'h0007E000;
                                              char44_2[38] <= 32'h0007E000;
                                              char44_2[39] <= 32'h0007E000;
                                              char44_2[40] <= 32'h0007E000;
                                              char44_2[41] <= 32'h0007E000;
                                              char44_2[42] <= 32'h0007E000;
                                              char44_2[43] <= 32'h0007E000;
                                              char44_2[44] <= 32'h0007E000;
                                              char44_2[45] <= 32'h0007E000;
                                              char44_2[46] <= 32'h0007E000;
                                              char44_2[47] <= 32'h0007E000;
                                              char44_2[48] <= 32'h0007E000;
                                              char44_2[49] <= 32'h0007E000;
                                              char44_2[50] <= 32'h0007E000;
                                              char44_2[51] <= 32'h000FF800;
                                              char44_2[52] <= 32'h03FFFFC0;
                                              char44_2[53] <= 32'h03FFFFC0;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//1
                                          4'd2: begin
                                              char44_2[  0] <= 32'h00000000;
                                              char44_2[  1] <= 32'h00000000;
                                              char44_2[  2] <= 32'h00000000;
                                              char44_2[  3] <= 32'h00000000;
                                              char44_2[  4] <= 32'h00000000;
                                              char44_2[  5] <= 32'h00000000;
                                              char44_2[  6] <= 32'h00000000;
                                              char44_2[  7] <= 32'h00000000;
                                              char44_2[  8] <= 32'h00000000;
                                              char44_2[  9] <= 32'h00000000;
                                              char44_2[10] <= 32'h001FFC00;
                                              char44_2[11] <= 32'h007FFF00;
                                              char44_2[12] <= 32'h01F83F80;
                                              char44_2[13] <= 32'h03E00FC0;
                                              char44_2[14] <= 32'h07C007E0;
                                              char44_2[15] <= 32'h078007E0;
                                              char44_2[16] <= 32'h0F8003F0;
                                              char44_2[17] <= 32'h0F8003F0;
                                              char44_2[18] <= 32'h1F8003F0;
                                              char44_2[19] <= 32'h1F8003F0;
                                              char44_2[20] <= 32'h1FC003F0;
                                              char44_2[21] <= 32'h1FC003F0;
                                              char44_2[22] <= 32'h1FC003F0;
                                              char44_2[23] <= 32'h0FC003F0;
                                              char44_2[24] <= 32'h07C003F0;
                                              char44_2[25] <= 32'h000003E0;
                                              char44_2[26] <= 32'h000007E0;
                                              char44_2[27] <= 32'h000007E0;
                                              char44_2[28] <= 32'h00000FC0;
                                              char44_2[29] <= 32'h00000F80;
                                              char44_2[30] <= 32'h00001F80;
                                              char44_2[31] <= 32'h00003F00;
                                              char44_2[32] <= 32'h00003E00;
                                              char44_2[33] <= 32'h00007C00;
                                              char44_2[34] <= 32'h0000F800;
                                              char44_2[35] <= 32'h0001F000;
                                              char44_2[36] <= 32'h0003E000;
                                              char44_2[37] <= 32'h0007C000;
                                              char44_2[38] <= 32'h000F8000;
                                              char44_2[39] <= 32'h001F0000;
                                              char44_2[40] <= 32'h003E0000;
                                              char44_2[41] <= 32'h007C0000;
                                              char44_2[42] <= 32'h00F80000;
                                              char44_2[43] <= 32'h01F00038;
                                              char44_2[44] <= 32'h01E00038;
                                              char44_2[45] <= 32'h03C00070;
                                              char44_2[46] <= 32'h07800070;
                                              char44_2[47] <= 32'h0F8000F0;
                                              char44_2[48] <= 32'h0F0000F0;
                                              char44_2[49] <= 32'h1E0003F0;
                                              char44_2[50] <= 32'h3FFFFFF0;
                                              char44_2[51] <= 32'h3FFFFFF0;
                                              char44_2[52] <= 32'h3FFFFFE0;
                                              char44_2[53] <= 32'h3FFFFFE0;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//2
                                          4'd3: begin
                                              char44_2[  0] <= 32'h00000000;
                                              char44_2[  1] <= 32'h00000000;
                                              char44_2[  2] <= 32'h00000000;
                                              char44_2[  3] <= 32'h00000000;
                                              char44_2[  4] <= 32'h00000000;
                                              char44_2[  5] <= 32'h00000000;
                                              char44_2[  6] <= 32'h00000000;
                                              char44_2[  7] <= 32'h00000000;
                                              char44_2[  8] <= 32'h00000000;
                                              char44_2[  9] <= 32'h00000000;
                                              char44_2[10] <= 32'h003FF000;
                                              char44_2[11] <= 32'h00FFFC00;
                                              char44_2[12] <= 32'h01F07E00;
                                              char44_2[13] <= 32'h03C03F00;
                                              char44_2[14] <= 32'h07801F80;
                                              char44_2[15] <= 32'h0F800FC0;
                                              char44_2[16] <= 32'h0F800FC0;
                                              char44_2[17] <= 32'h0F8007E0;
                                              char44_2[18] <= 32'h0FC007E0;
                                              char44_2[19] <= 32'h0FC007E0;
                                              char44_2[20] <= 32'h0FC007E0;
                                              char44_2[21] <= 32'h07C007E0;
                                              char44_2[22] <= 32'h000007E0;
                                              char44_2[23] <= 32'h000007E0;
                                              char44_2[24] <= 32'h000007C0;
                                              char44_2[25] <= 32'h00000FC0;
                                              char44_2[26] <= 32'h00000F80;
                                              char44_2[27] <= 32'h00001F00;
                                              char44_2[28] <= 32'h00007E00;
                                              char44_2[29] <= 32'h0003FC00;
                                              char44_2[30] <= 32'h001FF000;
                                              char44_2[31] <= 32'h001FFC00;
                                              char44_2[32] <= 32'h0000FF00;
                                              char44_2[33] <= 32'h00001F80;
                                              char44_2[34] <= 32'h00000FC0;
                                              char44_2[35] <= 32'h000007E0;
                                              char44_2[36] <= 32'h000003E0;
                                              char44_2[37] <= 32'h000003F0;
                                              char44_2[38] <= 32'h000003F0;
                                              char44_2[39] <= 32'h000001F0;
                                              char44_2[40] <= 32'h000001F8;
                                              char44_2[41] <= 32'h000001F8;
                                              char44_2[42] <= 32'h078001F8;
                                              char44_2[43] <= 32'h0FC001F8;
                                              char44_2[44] <= 32'h1FC001F8;
                                              char44_2[45] <= 32'h1FC003F0;
                                              char44_2[46] <= 32'h1FC003F0;
                                              char44_2[47] <= 32'h1FC003E0;
                                              char44_2[48] <= 32'h0F8007E0;
                                              char44_2[49] <= 32'h0F8007C0;
                                              char44_2[50] <= 32'h07C01F80;
                                              char44_2[51] <= 32'h03F07F00;
                                              char44_2[52] <= 32'h01FFFE00;
                                              char44_2[53] <= 32'h003FF000;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//3
                                          4'd4: begin
                                              char44_2[  0] <= 32'h00000000;
                                              char44_2[  1] <= 32'h00000000;
                                              char44_2[  2] <= 32'h00000000;
                                              char44_2[  3] <= 32'h00000000;
                                              char44_2[  4] <= 32'h00000000;
                                              char44_2[  5] <= 32'h00000000;
                                              char44_2[  6] <= 32'h00000000;
                                              char44_2[  7] <= 32'h00000000;
                                              char44_2[  8] <= 32'h00000000;
                                              char44_2[  9] <= 32'h00000000;
                                              char44_2[10] <= 32'h00001F00;
                                              char44_2[11] <= 32'h00001F00;
                                              char44_2[12] <= 32'h00003F00;
                                              char44_2[13] <= 32'h00003F00;
                                              char44_2[14] <= 32'h00007F00;
                                              char44_2[15] <= 32'h0000FF00;
                                              char44_2[16] <= 32'h0000FF00;
                                              char44_2[17] <= 32'h0001FF00;
                                              char44_2[18] <= 32'h0003FF00;
                                              char44_2[19] <= 32'h0003BF00;
                                              char44_2[20] <= 32'h0007BF00;
                                              char44_2[21] <= 32'h00073F00;
                                              char44_2[22] <= 32'h000F3F00;
                                              char44_2[23] <= 32'h001E3F00;
                                              char44_2[24] <= 32'h001C3F00;
                                              char44_2[25] <= 32'h003C3F00;
                                              char44_2[26] <= 32'h00783F00;
                                              char44_2[27] <= 32'h00783F00;
                                              char44_2[28] <= 32'h00F03F00;
                                              char44_2[29] <= 32'h00E03F00;
                                              char44_2[30] <= 32'h01E03F00;
                                              char44_2[31] <= 32'h03C03F00;
                                              char44_2[32] <= 32'h03803F00;
                                              char44_2[33] <= 32'h07803F00;
                                              char44_2[34] <= 32'h0F003F00;
                                              char44_2[35] <= 32'h0F003F00;
                                              char44_2[36] <= 32'h1E003F00;
                                              char44_2[37] <= 32'h1C003F00;
                                              char44_2[38] <= 32'h3C003F00;
                                              char44_2[39] <= 32'h7FFFFFFE;
                                              char44_2[40] <= 32'h7FFFFFFE;
                                              char44_2[41] <= 32'h00003F00;
                                              char44_2[42] <= 32'h00003F00;
                                              char44_2[43] <= 32'h00003F00;
                                              char44_2[44] <= 32'h00003F00;
                                              char44_2[45] <= 32'h00003F00;
                                              char44_2[46] <= 32'h00003F00;
                                              char44_2[47] <= 32'h00003F00;
                                              char44_2[48] <= 32'h00003F00;
                                              char44_2[49] <= 32'h00003F00;
                                              char44_2[50] <= 32'h00003F00;
                                              char44_2[51] <= 32'h00007F80;
                                              char44_2[52] <= 32'h000FFFFC;
                                              char44_2[53] <= 32'h000FFFFC;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//4
                                          4'd5: begin
                                              char44_2[  0] <= 32'h00000000;
                                              char44_2[  1] <= 32'h00000000;
                                              char44_2[  2] <= 32'h00000000;
                                              char44_2[  3] <= 32'h00000000;
                                              char44_2[  4] <= 32'h00000000;
                                              char44_2[  5] <= 32'h00000000;
                                              char44_2[  6] <= 32'h00000000;
                                              char44_2[  7] <= 32'h00000000;
                                              char44_2[  8] <= 32'h00000000;
                                              char44_2[  9] <= 32'h00000000;
                                              char44_2[10] <= 32'h00000000;
                                              char44_2[11] <= 32'h03FFFFF0;
                                              char44_2[12] <= 32'h03FFFFF0;
                                              char44_2[13] <= 32'h03FFFFF0;
                                              char44_2[14] <= 32'h03FFFFE0;
                                              char44_2[15] <= 32'h03800000;
                                              char44_2[16] <= 32'h03800000;
                                              char44_2[17] <= 32'h03800000;
                                              char44_2[18] <= 32'h03800000;
                                              char44_2[19] <= 32'h03800000;
                                              char44_2[20] <= 32'h07800000;
                                              char44_2[21] <= 32'h07800000;
                                              char44_2[22] <= 32'h07800000;
                                              char44_2[23] <= 32'h07800000;
                                              char44_2[24] <= 32'h07800000;
                                              char44_2[25] <= 32'h07800000;
                                              char44_2[26] <= 32'h078FF800;
                                              char44_2[27] <= 32'h073FFE00;
                                              char44_2[28] <= 32'h077FFF80;
                                              char44_2[29] <= 32'h07FC3F80;
                                              char44_2[30] <= 32'h07E00FC0;
                                              char44_2[31] <= 32'h07C007E0;
                                              char44_2[32] <= 32'h078007E0;
                                              char44_2[33] <= 32'h078003F0;
                                              char44_2[34] <= 32'h000003F0;
                                              char44_2[35] <= 32'h000001F0;
                                              char44_2[36] <= 32'h000001F8;
                                              char44_2[37] <= 32'h000001F8;
                                              char44_2[38] <= 32'h000001F8;
                                              char44_2[39] <= 32'h000001F8;
                                              char44_2[40] <= 32'h000001F8;
                                              char44_2[41] <= 32'h078001F8;
                                              char44_2[42] <= 32'h0FC001F8;
                                              char44_2[43] <= 32'h1FC001F0;
                                              char44_2[44] <= 32'h1FC001F0;
                                              char44_2[45] <= 32'h1FC003F0;
                                              char44_2[46] <= 32'h1F8003F0;
                                              char44_2[47] <= 32'h1F8003E0;
                                              char44_2[48] <= 32'h0F8007E0;
                                              char44_2[49] <= 32'h078007C0;
                                              char44_2[50] <= 32'h07C01F80;
                                              char44_2[51] <= 32'h03F83F00;
                                              char44_2[52] <= 32'h00FFFE00;
                                              char44_2[53] <= 32'h003FF800;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//5
                                          4'd6: begin
                                              char44_2[0] <= 32'h00000000;
                                              char44_2[1] <= 32'h00000000;
                                              char44_2[2] <= 32'h00000000;
                                              char44_2[3] <= 32'h00000000;
                                              char44_2[4] <= 32'h00000000;
                                              char44_2[5] <= 32'h00000000;
                                              char44_2[6] <= 32'h00000000;
                                              char44_2[7] <= 32'h00000000;
                                              char44_2[8] <= 32'h00000000;
                                              char44_2[9] <= 32'h00000000;
                                              char44_2[10] <= 32'h0007FE00;
                                              char44_2[11] <= 32'h001FFF80;
                                              char44_2[12] <= 32'h003F0FC0;
                                              char44_2[13] <= 32'h007C07C0;
                                              char44_2[14] <= 32'h00F807E0;
                                              char44_2[15] <= 32'h01F007E0;
                                              char44_2[16] <= 32'h03E007E0;
                                              char44_2[17] <= 32'h03C007E0;
                                              char44_2[18] <= 32'h07C003C0;
                                              char44_2[19] <= 32'h07C00000;
                                              char44_2[20] <= 32'h0FC00000;
                                              char44_2[21] <= 32'h0F800000;
                                              char44_2[22] <= 32'h0F800000;
                                              char44_2[23] <= 32'h1F800000;
                                              char44_2[24] <= 32'h1F800000;
                                              char44_2[25] <= 32'h1F800000;
                                              char44_2[26] <= 32'h1F87FE00;
                                              char44_2[27] <= 32'h1F9FFF80;
                                              char44_2[28] <= 32'h1FBFFFC0;
                                              char44_2[29] <= 32'h3FFE1FC0;
                                              char44_2[30] <= 32'h3FF807E0;
                                              char44_2[31] <= 32'h3FE003F0;
                                              char44_2[32] <= 32'h3FE003F0;
                                              char44_2[33] <= 32'h3FC001F8;
                                              char44_2[34] <= 32'h3F8001F8;
                                              char44_2[35] <= 32'h3F8001F8;
                                              char44_2[36] <= 32'h3F8000F8;
                                              char44_2[37] <= 32'h3F8000F8;
                                              char44_2[38] <= 32'h3F8000F8;
                                              char44_2[39] <= 32'h1F8000F8;
                                              char44_2[40] <= 32'h1F8000F8;
                                              char44_2[41] <= 32'h1F8000F8;
                                              char44_2[42] <= 32'h1F8000F8;
                                              char44_2[43] <= 32'h1F8000F8;
                                              char44_2[44] <= 32'h0FC001F8;
                                              char44_2[45] <= 32'h0FC001F8;
                                              char44_2[46] <= 32'h0FC001F0;
                                              char44_2[47] <= 32'h07E001F0;
                                              char44_2[48] <= 32'h03E003E0;
                                              char44_2[49] <= 32'h03F003E0;
                                              char44_2[50] <= 32'h01F807C0;
                                              char44_2[51] <= 32'h00FE1F80;
                                              char44_2[52] <= 32'h007FFE00;
                                              char44_2[53] <= 32'h001FF800;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//6
                                          4'd7: begin
                                              char44_2[0] <= 32'h00000000;
                                              char44_2[1] <= 32'h00000000;
                                              char44_2[2] <= 32'h00000000;
                                              char44_2[3] <= 32'h00000000;
                                              char44_2[4] <= 32'h00000000;
                                              char44_2[5] <= 32'h00000000;
                                              char44_2[6] <= 32'h00000000;
                                              char44_2[7] <= 32'h00000000;
                                              char44_2[8] <= 32'h00000000;
                                              char44_2[9] <= 32'h00000000;
                                              char44_2[10] <= 32'h00000000;
                                              char44_2[11] <= 32'h07FFFFF8;
                                              char44_2[12] <= 32'h07FFFFF8;
                                              char44_2[13] <= 32'h07FFFFF8;
                                              char44_2[14] <= 32'h0FFFFFF0;
                                              char44_2[15] <= 32'h0FC000E0;
                                              char44_2[16] <= 32'h0F8001E0;
                                              char44_2[17] <= 32'h0F0001C0;
                                              char44_2[18] <= 32'h0E0003C0;
                                              char44_2[19] <= 32'h0E000780;
                                              char44_2[20] <= 32'h1E000780;
                                              char44_2[21] <= 32'h1C000F00;
                                              char44_2[22] <= 32'h00000F00;
                                              char44_2[23] <= 32'h00001E00;
                                              char44_2[24] <= 32'h00001E00;
                                              char44_2[25] <= 32'h00003C00;
                                              char44_2[26] <= 32'h00003C00;
                                              char44_2[27] <= 32'h00007800;
                                              char44_2[28] <= 32'h00007800;
                                              char44_2[29] <= 32'h0000F800;
                                              char44_2[30] <= 32'h0000F000;
                                              char44_2[31] <= 32'h0001F000;
                                              char44_2[32] <= 32'h0001E000;
                                              char44_2[33] <= 32'h0003E000;
                                              char44_2[34] <= 32'h0003E000;
                                              char44_2[35] <= 32'h0003E000;
                                              char44_2[36] <= 32'h0007C000;
                                              char44_2[37] <= 32'h0007C000;
                                              char44_2[38] <= 32'h0007C000;
                                              char44_2[39] <= 32'h000FC000;
                                              char44_2[40] <= 32'h000FC000;
                                              char44_2[41] <= 32'h000FC000;
                                              char44_2[42] <= 32'h000FC000;
                                              char44_2[43] <= 32'h001FC000;
                                              char44_2[44] <= 32'h001FC000;
                                              char44_2[45] <= 32'h001FC000;
                                              char44_2[46] <= 32'h001FC000;
                                              char44_2[47] <= 32'h001FC000;
                                              char44_2[48] <= 32'h001FC000;
                                              char44_2[49] <= 32'h001FC000;
                                              char44_2[50] <= 32'h001FC000;
                                              char44_2[51] <= 32'h001FC000;
                                              char44_2[52] <= 32'h001FC000;
                                              char44_2[53] <= 32'h000F8000;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//7
                                          4'd8: begin
                                              char44_2[0] <= 32'h00000000;
                                              char44_2[1] <= 32'h00000000;
                                              char44_2[2] <= 32'h00000000;
                                              char44_2[3] <= 32'h00000000;
                                              char44_2[4] <= 32'h00000000;
                                              char44_2[5] <= 32'h00000000;
                                              char44_2[6] <= 32'h00000000;
                                              char44_2[7] <= 32'h00000000;
                                              char44_2[8] <= 32'h00000000;
                                              char44_2[9] <= 32'h00000000;
                                              char44_2[10] <= 32'h003FF800;
                                              char44_2[11] <= 32'h00FFFE00;
                                              char44_2[12] <= 32'h01F81F80;
                                              char44_2[13] <= 32'h03E00FC0;
                                              char44_2[14] <= 32'h07C003E0;
                                              char44_2[15] <= 32'h0F8003E0;
                                              char44_2[16] <= 32'h0F8001F0;
                                              char44_2[17] <= 32'h1F0001F0;
                                              char44_2[18] <= 32'h1F0001F0;
                                              char44_2[19] <= 32'h1F0001F0;
                                              char44_2[20] <= 32'h1F0001F0;
                                              char44_2[21] <= 32'h1F0001F0;
                                              char44_2[22] <= 32'h1F8001F0;
                                              char44_2[23] <= 32'h1FC001F0;
                                              char44_2[24] <= 32'h0FC001F0;
                                              char44_2[25] <= 32'h0FF003E0;
                                              char44_2[26] <= 32'h07F803C0;
                                              char44_2[27] <= 32'h03FE0F80;
                                              char44_2[28] <= 32'h01FF9F00;
                                              char44_2[29] <= 32'h00FFFE00;
                                              char44_2[30] <= 32'h003FF800;
                                              char44_2[31] <= 32'h007FFC00;
                                              char44_2[32] <= 32'h01F7FF00;
                                              char44_2[33] <= 32'h03E1FF80;
                                              char44_2[34] <= 32'h07C07FC0;
                                              char44_2[35] <= 32'h0F801FE0;
                                              char44_2[36] <= 32'h0F800FE0;
                                              char44_2[37] <= 32'h1F0007F0;
                                              char44_2[38] <= 32'h1F0003F0;
                                              char44_2[39] <= 32'h3E0001F8;
                                              char44_2[40] <= 32'h3E0001F8;
                                              char44_2[41] <= 32'h3E0001F8;
                                              char44_2[42] <= 32'h3E0000F8;
                                              char44_2[43] <= 32'h3E0000F8;
                                              char44_2[44] <= 32'h3E0000F8;
                                              char44_2[45] <= 32'h3E0000F8;
                                              char44_2[46] <= 32'h1F0001F0;
                                              char44_2[47] <= 32'h1F0001F0;
                                              char44_2[48] <= 32'h0F8003E0;
                                              char44_2[49] <= 32'h0FC003E0;
                                              char44_2[50] <= 32'h07E007C0;
                                              char44_2[51] <= 32'h01F83F80;
                                              char44_2[52] <= 32'h00FFFE00;
                                              char44_2[53] <= 32'h003FF800;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//8
                                          4'd9: begin
                                              char44_2[0] <= 32'h00000000;
                                              char44_2[1] <= 32'h00000000;
                                              char44_2[2] <= 32'h00000000;
                                              char44_2[3] <= 32'h00000000;
                                              char44_2[4] <= 32'h00000000;
                                              char44_2[5] <= 32'h00000000;
                                              char44_2[6] <= 32'h00000000;
                                              char44_2[7] <= 32'h00000000;
                                              char44_2[8] <= 32'h00000000;
                                              char44_2[9] <= 32'h00000000;
                                              char44_2[10] <= 32'h003FF000;
                                              char44_2[11] <= 32'h00FFFC00;
                                              char44_2[12] <= 32'h01F83F00;
                                              char44_2[13] <= 32'h03E01F80;
                                              char44_2[14] <= 32'h07C00F80;
                                              char44_2[15] <= 32'h0FC007C0;
                                              char44_2[16] <= 32'h0F8003E0;
                                              char44_2[17] <= 32'h1F8003E0;
                                              char44_2[18] <= 32'h1F0003F0;
                                              char44_2[19] <= 32'h1F0003F0;
                                              char44_2[20] <= 32'h3F0001F0;
                                              char44_2[21] <= 32'h3F0001F0;
                                              char44_2[22] <= 32'h3F0001F8;
                                              char44_2[23] <= 32'h3F0001F8;
                                              char44_2[24] <= 32'h3F0001F8;
                                              char44_2[25] <= 32'h3F0001F8;
                                              char44_2[26] <= 32'h3F0001F8;
                                              char44_2[27] <= 32'h3F0001F8;
                                              char44_2[28] <= 32'h3F0003F8;
                                              char44_2[29] <= 32'h1F8003F8;
                                              char44_2[30] <= 32'h1F8007F8;
                                              char44_2[31] <= 32'h1F800FF8;
                                              char44_2[32] <= 32'h0FC01FF8;
                                              char44_2[33] <= 32'h0FE03FF8;
                                              char44_2[34] <= 32'h07F8FDF8;
                                              char44_2[35] <= 32'h03FFF9F8;
                                              char44_2[36] <= 32'h01FFF1F8;
                                              char44_2[37] <= 32'h003F83F8;
                                              char44_2[38] <= 32'h000003F0;
                                              char44_2[39] <= 32'h000003F0;
                                              char44_2[40] <= 32'h000003F0;
                                              char44_2[41] <= 32'h000003F0;
                                              char44_2[42] <= 32'h000007E0;
                                              char44_2[43] <= 32'h000007E0;
                                              char44_2[44] <= 32'h000007C0;
                                              char44_2[45] <= 32'h03C007C0;
                                              char44_2[46] <= 32'h07C00F80;
                                              char44_2[47] <= 32'h0FE00F80;
                                              char44_2[48] <= 32'h0FE01F00;
                                              char44_2[49] <= 32'h0FE03E00;
                                              char44_2[50] <= 32'h07E07E00;
                                              char44_2[51] <= 32'h07F1F800;
                                              char44_2[52] <= 32'h03FFF000;
                                              char44_2[53] <= 32'h00FFC000;
                                              char44_2[54] <= 32'h00000000;
                                              char44_2[55] <= 32'h00000000;
                                              char44_2[56] <= 32'h00000000;
                                              char44_2[57] <= 32'h00000000;
                                              char44_2[58] <= 32'h00000000;
                                              char44_2[59] <= 32'h00000000;
                                              char44_2[60] <= 32'h00000000;
                                              char44_2[61] <= 32'h00000000;
                                              char44_2[62] <= 32'h00000000;
                                              char44_2[63] <= 32'h00000000;
                                          end//9
                                          default: begin
                                              char44_2[0] <= char44_2[0];
                                              char44_2[1] <= char44_2[1];
                                              char44_2[2] <= char44_2[2];
                                              char44_2[3] <= char44_2[3];
                                              char44_2[4] <= char44_2[4];
                                              char44_2[5] <= char44_2[5];
                                              char44_2[6] <= char44_2[6];
                                              char44_2[7] <= char44_2[7];
                                              char44_2[8] <= char44_2[8];
                                              char44_2[9] <= char44_2[9];
                                              char44_2[10] <= char44_2[10];
                                              char44_2[11] <= char44_2[11];
                                              char44_2[12] <= char44_2[12];
                                              char44_2[13] <= char44_2[13];
                                              char44_2[14] <= char44_2[14];
                                              char44_2[15] <= char44_2[15];
                                              char44_2[16] <= char44_2[16];
                                              char44_2[17] <= char44_2[17];
                                              char44_2[18] <= char44_2[18];
                                              char44_2[19] <= char44_2[19];
                                              char44_2[20] <= char44_2[20];
                                              char44_2[21] <= char44_2[21];
                                              char44_2[22] <= char44_2[22];
                                              char44_2[23] <= char44_2[23];
                                              char44_2[24] <= char44_2[24];
                                              char44_2[25] <= char44_2[25];
                                              char44_2[26] <= char44_2[26];
                                              char44_2[27] <= char44_2[27];
                                              char44_2[28] <= char44_2[28];
                                              char44_2[29] <= char44_2[29];
                                              char44_2[30] <= char44_2[30];
                                              char44_2[31] <= char44_2[31];
                                              char44_2[32] <= char44_2[32];
                                              char44_2[33] <= char44_2[33];
                                              char44_2[34] <= char44_2[34];
                                              char44_2[35] <= char44_2[35];
                                              char44_2[36] <= char44_2[36];
                                              char44_2[37] <= char44_2[37];
                                              char44_2[38] <= char44_2[38];
                                              char44_2[39] <= char44_2[39];
                                              char44_2[40] <= char44_2[40];
                                              char44_2[41] <= char44_2[41];
                                              char44_2[42] <= char44_2[42];
                                              char44_2[43] <= char44_2[43];
                                              char44_2[44] <= char44_2[44];
                                              char44_2[45] <= char44_2[45];
                                              char44_2[46] <= char44_2[46];
                                              char44_2[47] <= char44_2[47];
                                              char44_2[48] <= char44_2[48];
                                              char44_2[49] <= char44_2[49];
                                              char44_2[50] <= char44_2[50];
                                              char44_2[51] <= char44_2[51];
                                              char44_2[52] <= char44_2[52];
                                              char44_2[53] <= char44_2[53];
                                              char44_2[54] <= char44_2[54];
                                              char44_2[55] <= char44_2[55];
                                              char44_2[56] <= char44_2[56];
                                              char44_2[57] <= char44_2[57];
                                              char44_2[58] <= char44_2[58];
                                              char44_2[59] <= char44_2[59];
                                              char44_2[60] <= char44_2[60];
                                              char44_2[61] <= char44_2[61];
                                              char44_2[62] <= char44_2[62];
                                              char44_2[63] <= char44_2[63];
                                          end
                                      endcase
                          
                               case((a2 - h1*(a2/h1))/t1)
                                              4'd0: begin
                                                  char44_3[  0] <= 32'h00000000;
                                                  char44_3[  1] <= 32'h00000000;
                                                  char44_3[  2] <= 32'h00000000;
                                                  char44_3[  3] <= 32'h00000000;
                                                  char44_3[  4] <= 32'h00000000;
                                                  char44_3[  5] <= 32'h00000000;
                                                  char44_3[  6] <= 32'h00000000;
                                                  char44_3[  7] <= 32'h00000000;
                                                  char44_3[  8] <= 32'h00000000;
                                                  char44_3[  9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h000FF000;
                                                  char44_3[11] <= 32'h003FFC00;
                                                  char44_3[12] <= 32'h007E7E00;
                                                  char44_3[13] <= 32'h00F81F00;
                                                  char44_3[14] <= 32'h01F00F80;
                                                  char44_3[15] <= 32'h03F00FC0;
                                                  char44_3[16] <= 32'h03E007C0;
                                                  char44_3[17] <= 32'h07E007E0;
                                                  char44_3[18] <= 32'h07C003E0;
                                                  char44_3[19] <= 32'h0FC003F0;
                                                  char44_3[20] <= 32'h0FC003F0;
                                                  char44_3[21] <= 32'h0FC003F0;
                                                  char44_3[22] <= 32'h1F8001F8;
                                                  char44_3[23] <= 32'h1F8001F8;
                                                  char44_3[24] <= 32'h1F8001F8;
                                                  char44_3[25] <= 32'h1F8001F8;
                                                  char44_3[26] <= 32'h1F8001F8;
                                                  char44_3[27] <= 32'h3F8001F8;
                                                  char44_3[28] <= 32'h3F8001F8;
                                                  char44_3[29] <= 32'h3F8001F8;
                                                  char44_3[30] <= 32'h3F8001F8;
                                                  char44_3[31] <= 32'h3F8001F8;
                                                  char44_3[32] <= 32'h3F8001F8;
                                                  char44_3[33] <= 32'h3F8001F8;
                                                  char44_3[34] <= 32'h3F8001F8;
                                                  char44_3[35] <= 32'h3F8001F8;
                                                  char44_3[36] <= 32'h3F8001F8;
                                                  char44_3[37] <= 32'h1F8001F8;
                                                  char44_3[38] <= 32'h1F8001F8;
                                                  char44_3[39] <= 32'h1F8001F8;
                                                  char44_3[40] <= 32'h1F8001F8;
                                                  char44_3[41] <= 32'h1F8001F0;
                                                  char44_3[42] <= 32'h0F8003F0;
                                                  char44_3[43] <= 32'h0FC003F0;
                                                  char44_3[44] <= 32'h0FC003F0;
                                                  char44_3[45] <= 32'h07C003E0;
                                                  char44_3[46] <= 32'h07E007E0;
                                                  char44_3[47] <= 32'h03E007C0;
                                                  char44_3[48] <= 32'h03F00FC0;
                                                  char44_3[49] <= 32'h01F00F80;
                                                  char44_3[50] <= 32'h00F81F00;
                                                  char44_3[51] <= 32'h007E7E00;
                                                  char44_3[52] <= 32'h003FFC00;
                                                  char44_3[53] <= 32'h000FF000;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//0
                                              4'd1: begin
                                                  char44_3[  0] <= 32'h00000000;
                                                  char44_3[  1] <= 32'h00000000;
                                                  char44_3[  2] <= 32'h00000000;
                                                  char44_3[  3] <= 32'h00000000;
                                                  char44_3[  4] <= 32'h00000000;
                                                  char44_3[  5] <= 32'h00000000;
                                                  char44_3[  6] <= 32'h00000000;
                                                  char44_3[  7] <= 32'h00000000;
                                                  char44_3[  8] <= 32'h00000000;
                                                  char44_3[  9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h0000E000;
                                                  char44_3[11] <= 32'h0001E000;
                                                  char44_3[12] <= 32'h0003E000;
                                                  char44_3[13] <= 32'h001FE000;
                                                  char44_3[14] <= 32'h03FFE000;
                                                  char44_3[15] <= 32'h03FFE000;
                                                  char44_3[16] <= 32'h0007E000;
                                                  char44_3[17] <= 32'h0007E000;
                                                  char44_3[18] <= 32'h0007E000;
                                                  char44_3[19] <= 32'h0007E000;
                                                  char44_3[20] <= 32'h0007E000;
                                                  char44_3[21] <= 32'h0007E000;
                                                  char44_3[22] <= 32'h0007E000;
                                                  char44_3[23] <= 32'h0007E000;
                                                  char44_3[24] <= 32'h0007E000;
                                                  char44_3[25] <= 32'h0007E000;
                                                  char44_3[26] <= 32'h0007E000;
                                                  char44_3[27] <= 32'h0007E000;
                                                  char44_3[28] <= 32'h0007E000;
                                                  char44_3[29] <= 32'h0007E000;
                                                  char44_3[30] <= 32'h0007E000;
                                                  char44_3[31] <= 32'h0007E000;
                                                  char44_3[32] <= 32'h0007E000;
                                                  char44_3[33] <= 32'h0007E000;
                                                  char44_3[34] <= 32'h0007E000;
                                                  char44_3[35] <= 32'h0007E000;
                                                  char44_3[36] <= 32'h0007E000;
                                                  char44_3[37] <= 32'h0007E000;
                                                  char44_3[38] <= 32'h0007E000;
                                                  char44_3[39] <= 32'h0007E000;
                                                  char44_3[40] <= 32'h0007E000;
                                                  char44_3[41] <= 32'h0007E000;
                                                  char44_3[42] <= 32'h0007E000;
                                                  char44_3[43] <= 32'h0007E000;
                                                  char44_3[44] <= 32'h0007E000;
                                                  char44_3[45] <= 32'h0007E000;
                                                  char44_3[46] <= 32'h0007E000;
                                                  char44_3[47] <= 32'h0007E000;
                                                  char44_3[48] <= 32'h0007E000;
                                                  char44_3[49] <= 32'h0007E000;
                                                  char44_3[50] <= 32'h0007E000;
                                                  char44_3[51] <= 32'h000FF800;
                                                  char44_3[52] <= 32'h03FFFFC0;
                                                  char44_3[53] <= 32'h03FFFFC0;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//1
                                              4'd2: begin
                                                  char44_3[  0] <= 32'h00000000;
                                                  char44_3[  1] <= 32'h00000000;
                                                  char44_3[  2] <= 32'h00000000;
                                                  char44_3[  3] <= 32'h00000000;
                                                  char44_3[  4] <= 32'h00000000;
                                                  char44_3[  5] <= 32'h00000000;
                                                  char44_3[  6] <= 32'h00000000;
                                                  char44_3[  7] <= 32'h00000000;
                                                  char44_3[  8] <= 32'h00000000;
                                                  char44_3[  9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h001FFC00;
                                                  char44_3[11] <= 32'h007FFF00;
                                                  char44_3[12] <= 32'h01F83F80;
                                                  char44_3[13] <= 32'h03E00FC0;
                                                  char44_3[14] <= 32'h07C007E0;
                                                  char44_3[15] <= 32'h078007E0;
                                                  char44_3[16] <= 32'h0F8003F0;
                                                  char44_3[17] <= 32'h0F8003F0;
                                                  char44_3[18] <= 32'h1F8003F0;
                                                  char44_3[19] <= 32'h1F8003F0;
                                                  char44_3[20] <= 32'h1FC003F0;
                                                  char44_3[21] <= 32'h1FC003F0;
                                                  char44_3[22] <= 32'h1FC003F0;
                                                  char44_3[23] <= 32'h0FC003F0;
                                                  char44_3[24] <= 32'h07C003F0;
                                                  char44_3[25] <= 32'h000003E0;
                                                  char44_3[26] <= 32'h000007E0;
                                                  char44_3[27] <= 32'h000007E0;
                                                  char44_3[28] <= 32'h00000FC0;
                                                  char44_3[29] <= 32'h00000F80;
                                                  char44_3[30] <= 32'h00001F80;
                                                  char44_3[31] <= 32'h00003F00;
                                                  char44_3[32] <= 32'h00003E00;
                                                  char44_3[33] <= 32'h00007C00;
                                                  char44_3[34] <= 32'h0000F800;
                                                  char44_3[35] <= 32'h0001F000;
                                                  char44_3[36] <= 32'h0003E000;
                                                  char44_3[37] <= 32'h0007C000;
                                                  char44_3[38] <= 32'h000F8000;
                                                  char44_3[39] <= 32'h001F0000;
                                                  char44_3[40] <= 32'h003E0000;
                                                  char44_3[41] <= 32'h007C0000;
                                                  char44_3[42] <= 32'h00F80000;
                                                  char44_3[43] <= 32'h01F00038;
                                                  char44_3[44] <= 32'h01E00038;
                                                  char44_3[45] <= 32'h03C00070;
                                                  char44_3[46] <= 32'h07800070;
                                                  char44_3[47] <= 32'h0F8000F0;
                                                  char44_3[48] <= 32'h0F0000F0;
                                                  char44_3[49] <= 32'h1E0003F0;
                                                  char44_3[50] <= 32'h3FFFFFF0;
                                                  char44_3[51] <= 32'h3FFFFFF0;
                                                  char44_3[52] <= 32'h3FFFFFE0;
                                                  char44_3[53] <= 32'h3FFFFFE0;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//2
                                              4'd3: begin
                                                  char44_3[  0] <= 32'h00000000;
                                                  char44_3[  1] <= 32'h00000000;
                                                  char44_3[  2] <= 32'h00000000;
                                                  char44_3[  3] <= 32'h00000000;
                                                  char44_3[  4] <= 32'h00000000;
                                                  char44_3[  5] <= 32'h00000000;
                                                  char44_3[  6] <= 32'h00000000;
                                                  char44_3[  7] <= 32'h00000000;
                                                  char44_3[  8] <= 32'h00000000;
                                                  char44_3[  9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h003FF000;
                                                  char44_3[11] <= 32'h00FFFC00;
                                                  char44_3[12] <= 32'h01F07E00;
                                                  char44_3[13] <= 32'h03C03F00;
                                                  char44_3[14] <= 32'h07801F80;
                                                  char44_3[15] <= 32'h0F800FC0;
                                                  char44_3[16] <= 32'h0F800FC0;
                                                  char44_3[17] <= 32'h0F8007E0;
                                                  char44_3[18] <= 32'h0FC007E0;
                                                  char44_3[19] <= 32'h0FC007E0;
                                                  char44_3[20] <= 32'h0FC007E0;
                                                  char44_3[21] <= 32'h07C007E0;
                                                  char44_3[22] <= 32'h000007E0;
                                                  char44_3[23] <= 32'h000007E0;
                                                  char44_3[24] <= 32'h000007C0;
                                                  char44_3[25] <= 32'h00000FC0;
                                                  char44_3[26] <= 32'h00000F80;
                                                  char44_3[27] <= 32'h00001F00;
                                                  char44_3[28] <= 32'h00007E00;
                                                  char44_3[29] <= 32'h0003FC00;
                                                  char44_3[30] <= 32'h001FF000;
                                                  char44_3[31] <= 32'h001FFC00;
                                                  char44_3[32] <= 32'h0000FF00;
                                                  char44_3[33] <= 32'h00001F80;
                                                  char44_3[34] <= 32'h00000FC0;
                                                  char44_3[35] <= 32'h000007E0;
                                                  char44_3[36] <= 32'h000003E0;
                                                  char44_3[37] <= 32'h000003F0;
                                                  char44_3[38] <= 32'h000003F0;
                                                  char44_3[39] <= 32'h000001F0;
                                                  char44_3[40] <= 32'h000001F8;
                                                  char44_3[41] <= 32'h000001F8;
                                                  char44_3[42] <= 32'h078001F8;
                                                  char44_3[43] <= 32'h0FC001F8;
                                                  char44_3[44] <= 32'h1FC001F8;
                                                  char44_3[45] <= 32'h1FC003F0;
                                                  char44_3[46] <= 32'h1FC003F0;
                                                  char44_3[47] <= 32'h1FC003E0;
                                                  char44_3[48] <= 32'h0F8007E0;
                                                  char44_3[49] <= 32'h0F8007C0;
                                                  char44_3[50] <= 32'h07C01F80;
                                                  char44_3[51] <= 32'h03F07F00;
                                                  char44_3[52] <= 32'h01FFFE00;
                                                  char44_3[53] <= 32'h003FF000;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//3
                                              4'd4: begin
                                                  char44_3[  0] <= 32'h00000000;
                                                  char44_3[  1] <= 32'h00000000;
                                                  char44_3[  2] <= 32'h00000000;
                                                  char44_3[  3] <= 32'h00000000;
                                                  char44_3[  4] <= 32'h00000000;
                                                  char44_3[  5] <= 32'h00000000;
                                                  char44_3[  6] <= 32'h00000000;
                                                  char44_3[  7] <= 32'h00000000;
                                                  char44_3[  8] <= 32'h00000000;
                                                  char44_3[  9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h00001F00;
                                                  char44_3[11] <= 32'h00001F00;
                                                  char44_3[12] <= 32'h00003F00;
                                                  char44_3[13] <= 32'h00003F00;
                                                  char44_3[14] <= 32'h00007F00;
                                                  char44_3[15] <= 32'h0000FF00;
                                                  char44_3[16] <= 32'h0000FF00;
                                                  char44_3[17] <= 32'h0001FF00;
                                                  char44_3[18] <= 32'h0003FF00;
                                                  char44_3[19] <= 32'h0003BF00;
                                                  char44_3[20] <= 32'h0007BF00;
                                                  char44_3[21] <= 32'h00073F00;
                                                  char44_3[22] <= 32'h000F3F00;
                                                  char44_3[23] <= 32'h001E3F00;
                                                  char44_3[24] <= 32'h001C3F00;
                                                  char44_3[25] <= 32'h003C3F00;
                                                  char44_3[26] <= 32'h00783F00;
                                                  char44_3[27] <= 32'h00783F00;
                                                  char44_3[28] <= 32'h00F03F00;
                                                  char44_3[29] <= 32'h00E03F00;
                                                  char44_3[30] <= 32'h01E03F00;
                                                  char44_3[31] <= 32'h03C03F00;
                                                  char44_3[32] <= 32'h03803F00;
                                                  char44_3[33] <= 32'h07803F00;
                                                  char44_3[34] <= 32'h0F003F00;
                                                  char44_3[35] <= 32'h0F003F00;
                                                  char44_3[36] <= 32'h1E003F00;
                                                  char44_3[37] <= 32'h1C003F00;
                                                  char44_3[38] <= 32'h3C003F00;
                                                  char44_3[39] <= 32'h7FFFFFFE;
                                                  char44_3[40] <= 32'h7FFFFFFE;
                                                  char44_3[41] <= 32'h00003F00;
                                                  char44_3[42] <= 32'h00003F00;
                                                  char44_3[43] <= 32'h00003F00;
                                                  char44_3[44] <= 32'h00003F00;
                                                  char44_3[45] <= 32'h00003F00;
                                                  char44_3[46] <= 32'h00003F00;
                                                  char44_3[47] <= 32'h00003F00;
                                                  char44_3[48] <= 32'h00003F00;
                                                  char44_3[49] <= 32'h00003F00;
                                                  char44_3[50] <= 32'h00003F00;
                                                  char44_3[51] <= 32'h00007F80;
                                                  char44_3[52] <= 32'h000FFFFC;
                                                  char44_3[53] <= 32'h000FFFFC;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//4
                                              4'd5: begin
                                                  char44_3[  0] <= 32'h00000000;
                                                  char44_3[  1] <= 32'h00000000;
                                                  char44_3[  2] <= 32'h00000000;
                                                  char44_3[  3] <= 32'h00000000;
                                                  char44_3[  4] <= 32'h00000000;
                                                  char44_3[  5] <= 32'h00000000;
                                                  char44_3[  6] <= 32'h00000000;
                                                  char44_3[  7] <= 32'h00000000;
                                                  char44_3[  8] <= 32'h00000000;
                                                  char44_3[  9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h00000000;
                                                  char44_3[11] <= 32'h03FFFFF0;
                                                  char44_3[12] <= 32'h03FFFFF0;
                                                  char44_3[13] <= 32'h03FFFFF0;
                                                  char44_3[14] <= 32'h03FFFFE0;
                                                  char44_3[15] <= 32'h03800000;
                                                  char44_3[16] <= 32'h03800000;
                                                  char44_3[17] <= 32'h03800000;
                                                  char44_3[18] <= 32'h03800000;
                                                  char44_3[19] <= 32'h03800000;
                                                  char44_3[20] <= 32'h07800000;
                                                  char44_3[21] <= 32'h07800000;
                                                  char44_3[22] <= 32'h07800000;
                                                  char44_3[23] <= 32'h07800000;
                                                  char44_3[24] <= 32'h07800000;
                                                  char44_3[25] <= 32'h07800000;
                                                  char44_3[26] <= 32'h078FF800;
                                                  char44_3[27] <= 32'h073FFE00;
                                                  char44_3[28] <= 32'h077FFF80;
                                                  char44_3[29] <= 32'h07FC3F80;
                                                  char44_3[30] <= 32'h07E00FC0;
                                                  char44_3[31] <= 32'h07C007E0;
                                                  char44_3[32] <= 32'h078007E0;
                                                  char44_3[33] <= 32'h078003F0;
                                                  char44_3[34] <= 32'h000003F0;
                                                  char44_3[35] <= 32'h000001F0;
                                                  char44_3[36] <= 32'h000001F8;
                                                  char44_3[37] <= 32'h000001F8;
                                                  char44_3[38] <= 32'h000001F8;
                                                  char44_3[39] <= 32'h000001F8;
                                                  char44_3[40] <= 32'h000001F8;
                                                  char44_3[41] <= 32'h078001F8;
                                                  char44_3[42] <= 32'h0FC001F8;
                                                  char44_3[43] <= 32'h1FC001F0;
                                                  char44_3[44] <= 32'h1FC001F0;
                                                  char44_3[45] <= 32'h1FC003F0;
                                                  char44_3[46] <= 32'h1F8003F0;
                                                  char44_3[47] <= 32'h1F8003E0;
                                                  char44_3[48] <= 32'h0F8007E0;
                                                  char44_3[49] <= 32'h078007C0;
                                                  char44_3[50] <= 32'h07C01F80;
                                                  char44_3[51] <= 32'h03F83F00;
                                                  char44_3[52] <= 32'h00FFFE00;
                                                  char44_3[53] <= 32'h003FF800;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//5
                                              4'd6: begin
                                                  char44_3[0] <= 32'h00000000;
                                                  char44_3[1] <= 32'h00000000;
                                                  char44_3[2] <= 32'h00000000;
                                                  char44_3[3] <= 32'h00000000;
                                                  char44_3[4] <= 32'h00000000;
                                                  char44_3[5] <= 32'h00000000;
                                                  char44_3[6] <= 32'h00000000;
                                                  char44_3[7] <= 32'h00000000;
                                                  char44_3[8] <= 32'h00000000;
                                                  char44_3[9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h0007FE00;
                                                  char44_3[11] <= 32'h001FFF80;
                                                  char44_3[12] <= 32'h003F0FC0;
                                                  char44_3[13] <= 32'h007C07C0;
                                                  char44_3[14] <= 32'h00F807E0;
                                                  char44_3[15] <= 32'h01F007E0;
                                                  char44_3[16] <= 32'h03E007E0;
                                                  char44_3[17] <= 32'h03C007E0;
                                                  char44_3[18] <= 32'h07C003C0;
                                                  char44_3[19] <= 32'h07C00000;
                                                  char44_3[20] <= 32'h0FC00000;
                                                  char44_3[21] <= 32'h0F800000;
                                                  char44_3[22] <= 32'h0F800000;
                                                  char44_3[23] <= 32'h1F800000;
                                                  char44_3[24] <= 32'h1F800000;
                                                  char44_3[25] <= 32'h1F800000;
                                                  char44_3[26] <= 32'h1F87FE00;
                                                  char44_3[27] <= 32'h1F9FFF80;
                                                  char44_3[28] <= 32'h1FBFFFC0;
                                                  char44_3[29] <= 32'h3FFE1FC0;
                                                  char44_3[30] <= 32'h3FF807E0;
                                                  char44_3[31] <= 32'h3FE003F0;
                                                  char44_3[32] <= 32'h3FE003F0;
                                                  char44_3[33] <= 32'h3FC001F8;
                                                  char44_3[34] <= 32'h3F8001F8;
                                                  char44_3[35] <= 32'h3F8001F8;
                                                  char44_3[36] <= 32'h3F8000F8;
                                                  char44_3[37] <= 32'h3F8000F8;
                                                  char44_3[38] <= 32'h3F8000F8;
                                                  char44_3[39] <= 32'h1F8000F8;
                                                  char44_3[40] <= 32'h1F8000F8;
                                                  char44_3[41] <= 32'h1F8000F8;
                                                  char44_3[42] <= 32'h1F8000F8;
                                                  char44_3[43] <= 32'h1F8000F8;
                                                  char44_3[44] <= 32'h0FC001F8;
                                                  char44_3[45] <= 32'h0FC001F8;
                                                  char44_3[46] <= 32'h0FC001F0;
                                                  char44_3[47] <= 32'h07E001F0;
                                                  char44_3[48] <= 32'h03E003E0;
                                                  char44_3[49] <= 32'h03F003E0;
                                                  char44_3[50] <= 32'h01F807C0;
                                                  char44_3[51] <= 32'h00FE1F80;
                                                  char44_3[52] <= 32'h007FFE00;
                                                  char44_3[53] <= 32'h001FF800;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//6
                                              4'd7: begin
                                                  char44_3[0] <= 32'h00000000;
                                                  char44_3[1] <= 32'h00000000;
                                                  char44_3[2] <= 32'h00000000;
                                                  char44_3[3] <= 32'h00000000;
                                                  char44_3[4] <= 32'h00000000;
                                                  char44_3[5] <= 32'h00000000;
                                                  char44_3[6] <= 32'h00000000;
                                                  char44_3[7] <= 32'h00000000;
                                                  char44_3[8] <= 32'h00000000;
                                                  char44_3[9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h00000000;
                                                  char44_3[11] <= 32'h07FFFFF8;
                                                  char44_3[12] <= 32'h07FFFFF8;
                                                  char44_3[13] <= 32'h07FFFFF8;
                                                  char44_3[14] <= 32'h0FFFFFF0;
                                                  char44_3[15] <= 32'h0FC000E0;
                                                  char44_3[16] <= 32'h0F8001E0;
                                                  char44_3[17] <= 32'h0F0001C0;
                                                  char44_3[18] <= 32'h0E0003C0;
                                                  char44_3[19] <= 32'h0E000780;
                                                  char44_3[20] <= 32'h1E000780;
                                                  char44_3[21] <= 32'h1C000F00;
                                                  char44_3[22] <= 32'h00000F00;
                                                  char44_3[23] <= 32'h00001E00;
                                                  char44_3[24] <= 32'h00001E00;
                                                  char44_3[25] <= 32'h00003C00;
                                                  char44_3[26] <= 32'h00003C00;
                                                  char44_3[27] <= 32'h00007800;
                                                  char44_3[28] <= 32'h00007800;
                                                  char44_3[29] <= 32'h0000F800;
                                                  char44_3[30] <= 32'h0000F000;
                                                  char44_3[31] <= 32'h0001F000;
                                                  char44_3[32] <= 32'h0001E000;
                                                  char44_3[33] <= 32'h0003E000;
                                                  char44_3[34] <= 32'h0003E000;
                                                  char44_3[35] <= 32'h0003E000;
                                                  char44_3[36] <= 32'h0007C000;
                                                  char44_3[37] <= 32'h0007C000;
                                                  char44_3[38] <= 32'h0007C000;
                                                  char44_3[39] <= 32'h000FC000;
                                                  char44_3[40] <= 32'h000FC000;
                                                  char44_3[41] <= 32'h000FC000;
                                                  char44_3[42] <= 32'h000FC000;
                                                  char44_3[43] <= 32'h001FC000;
                                                  char44_3[44] <= 32'h001FC000;
                                                  char44_3[45] <= 32'h001FC000;
                                                  char44_3[46] <= 32'h001FC000;
                                                  char44_3[47] <= 32'h001FC000;
                                                  char44_3[48] <= 32'h001FC000;
                                                  char44_3[49] <= 32'h001FC000;
                                                  char44_3[50] <= 32'h001FC000;
                                                  char44_3[51] <= 32'h001FC000;
                                                  char44_3[52] <= 32'h001FC000;
                                                  char44_3[53] <= 32'h000F8000;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//7
                                              4'd8: begin
                                                  char44_3[0] <= 32'h00000000;
                                                  char44_3[1] <= 32'h00000000;
                                                  char44_3[2] <= 32'h00000000;
                                                  char44_3[3] <= 32'h00000000;
                                                  char44_3[4] <= 32'h00000000;
                                                  char44_3[5] <= 32'h00000000;
                                                  char44_3[6] <= 32'h00000000;
                                                  char44_3[7] <= 32'h00000000;
                                                  char44_3[8] <= 32'h00000000;
                                                  char44_3[9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h003FF800;
                                                  char44_3[11] <= 32'h00FFFE00;
                                                  char44_3[12] <= 32'h01F81F80;
                                                  char44_3[13] <= 32'h03E00FC0;
                                                  char44_3[14] <= 32'h07C003E0;
                                                  char44_3[15] <= 32'h0F8003E0;
                                                  char44_3[16] <= 32'h0F8001F0;
                                                  char44_3[17] <= 32'h1F0001F0;
                                                  char44_3[18] <= 32'h1F0001F0;
                                                  char44_3[19] <= 32'h1F0001F0;
                                                  char44_3[20] <= 32'h1F0001F0;
                                                  char44_3[21] <= 32'h1F0001F0;
                                                  char44_3[22] <= 32'h1F8001F0;
                                                  char44_3[23] <= 32'h1FC001F0;
                                                  char44_3[24] <= 32'h0FC001F0;
                                                  char44_3[25] <= 32'h0FF003E0;
                                                  char44_3[26] <= 32'h07F803C0;
                                                  char44_3[27] <= 32'h03FE0F80;
                                                  char44_3[28] <= 32'h01FF9F00;
                                                  char44_3[29] <= 32'h00FFFE00;
                                                  char44_3[30] <= 32'h003FF800;
                                                  char44_3[31] <= 32'h007FFC00;
                                                  char44_3[32] <= 32'h01F7FF00;
                                                  char44_3[33] <= 32'h03E1FF80;
                                                  char44_3[34] <= 32'h07C07FC0;
                                                  char44_3[35] <= 32'h0F801FE0;
                                                  char44_3[36] <= 32'h0F800FE0;
                                                  char44_3[37] <= 32'h1F0007F0;
                                                  char44_3[38] <= 32'h1F0003F0;
                                                  char44_3[39] <= 32'h3E0001F8;
                                                  char44_3[40] <= 32'h3E0001F8;
                                                  char44_3[41] <= 32'h3E0001F8;
                                                  char44_3[42] <= 32'h3E0000F8;
                                                  char44_3[43] <= 32'h3E0000F8;
                                                  char44_3[44] <= 32'h3E0000F8;
                                                  char44_3[45] <= 32'h3E0000F8;
                                                  char44_3[46] <= 32'h1F0001F0;
                                                  char44_3[47] <= 32'h1F0001F0;
                                                  char44_3[48] <= 32'h0F8003E0;
                                                  char44_3[49] <= 32'h0FC003E0;
                                                  char44_3[50] <= 32'h07E007C0;
                                                  char44_3[51] <= 32'h01F83F80;
                                                  char44_3[52] <= 32'h00FFFE00;
                                                  char44_3[53] <= 32'h003FF800;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//8
                                              4'd9: begin
                                                  char44_3[0] <= 32'h00000000;
                                                  char44_3[1] <= 32'h00000000;
                                                  char44_3[2] <= 32'h00000000;
                                                  char44_3[3] <= 32'h00000000;
                                                  char44_3[4] <= 32'h00000000;
                                                  char44_3[5] <= 32'h00000000;
                                                  char44_3[6] <= 32'h00000000;
                                                  char44_3[7] <= 32'h00000000;
                                                  char44_3[8] <= 32'h00000000;
                                                  char44_3[9] <= 32'h00000000;
                                                  char44_3[10] <= 32'h003FF000;
                                                  char44_3[11] <= 32'h00FFFC00;
                                                  char44_3[12] <= 32'h01F83F00;
                                                  char44_3[13] <= 32'h03E01F80;
                                                  char44_3[14] <= 32'h07C00F80;
                                                  char44_3[15] <= 32'h0FC007C0;
                                                  char44_3[16] <= 32'h0F8003E0;
                                                  char44_3[17] <= 32'h1F8003E0;
                                                  char44_3[18] <= 32'h1F0003F0;
                                                  char44_3[19] <= 32'h1F0003F0;
                                                  char44_3[20] <= 32'h3F0001F0;
                                                  char44_3[21] <= 32'h3F0001F0;
                                                  char44_3[22] <= 32'h3F0001F8;
                                                  char44_3[23] <= 32'h3F0001F8;
                                                  char44_3[24] <= 32'h3F0001F8;
                                                  char44_3[25] <= 32'h3F0001F8;
                                                  char44_3[26] <= 32'h3F0001F8;
                                                  char44_3[27] <= 32'h3F0001F8;
                                                  char44_3[28] <= 32'h3F0003F8;
                                                  char44_3[29] <= 32'h1F8003F8;
                                                  char44_3[30] <= 32'h1F8007F8;
                                                  char44_3[31] <= 32'h1F800FF8;
                                                  char44_3[32] <= 32'h0FC01FF8;
                                                  char44_3[33] <= 32'h0FE03FF8;
                                                  char44_3[34] <= 32'h07F8FDF8;
                                                  char44_3[35] <= 32'h03FFF9F8;
                                                  char44_3[36] <= 32'h01FFF1F8;
                                                  char44_3[37] <= 32'h003F83F8;
                                                  char44_3[38] <= 32'h000003F0;
                                                  char44_3[39] <= 32'h000003F0;
                                                  char44_3[40] <= 32'h000003F0;
                                                  char44_3[41] <= 32'h000003F0;
                                                  char44_3[42] <= 32'h000007E0;
                                                  char44_3[43] <= 32'h000007E0;
                                                  char44_3[44] <= 32'h000007C0;
                                                  char44_3[45] <= 32'h03C007C0;
                                                  char44_3[46] <= 32'h07C00F80;
                                                  char44_3[47] <= 32'h0FE00F80;
                                                  char44_3[48] <= 32'h0FE01F00;
                                                  char44_3[49] <= 32'h0FE03E00;
                                                  char44_3[50] <= 32'h07E07E00;
                                                  char44_3[51] <= 32'h07F1F800;
                                                  char44_3[52] <= 32'h03FFF000;
                                                  char44_3[53] <= 32'h00FFC000;
                                                  char44_3[54] <= 32'h00000000;
                                                  char44_3[55] <= 32'h00000000;
                                                  char44_3[56] <= 32'h00000000;
                                                  char44_3[57] <= 32'h00000000;
                                                  char44_3[58] <= 32'h00000000;
                                                  char44_3[59] <= 32'h00000000;
                                                  char44_3[60] <= 32'h00000000;
                                                  char44_3[61] <= 32'h00000000;
                                                  char44_3[62] <= 32'h00000000;
                                                  char44_3[63] <= 32'h00000000;
                                              end//9
                                              default: begin
                                                  char44_3[0] <= char44_3[0];
                                                  char44_3[1] <= char44_3[1];
                                                  char44_3[2] <= char44_3[2];
                                                  char44_3[3] <= char44_3[3];
                                                  char44_3[4] <= char44_3[4];
                                                  char44_3[5] <= char44_3[5];
                                                  char44_3[6] <= char44_3[6];
                                                  char44_3[7] <= char44_3[7];
                                                  char44_3[8] <= char44_3[8];
                                                  char44_3[9] <= char44_3[9];
                                                  char44_3[10] <= char44_3[10];
                                                  char44_3[11] <= char44_3[11];
                                                  char44_3[12] <= char44_3[12];
                                                  char44_3[13] <= char44_3[13];
                                                  char44_3[14] <= char44_3[14];
                                                  char44_3[15] <= char44_3[15];
                                                  char44_3[16] <= char44_3[16];
                                                  char44_3[17] <= char44_3[17];
                                                  char44_3[18] <= char44_3[18];
                                                  char44_3[19] <= char44_3[19];
                                                  char44_3[20] <= char44_3[20];
                                                  char44_3[21] <= char44_3[21];
                                                  char44_3[22] <= char44_3[22];
                                                  char44_3[23] <= char44_3[23];
                                                  char44_3[24] <= char44_3[24];
                                                  char44_3[25] <= char44_3[25];
                                                  char44_3[26] <= char44_3[26];
                                                  char44_3[27] <= char44_3[27];
                                                  char44_3[28] <= char44_3[28];
                                                  char44_3[29] <= char44_3[29];
                                                  char44_3[30] <= char44_3[30];
                                                  char44_3[31] <= char44_3[31];
                                                  char44_3[32] <= char44_3[32];
                                                  char44_3[33] <= char44_3[33];
                                                  char44_3[34] <= char44_3[34];
                                                  char44_3[35] <= char44_3[35];
                                                  char44_3[36] <= char44_3[36];
                                                  char44_3[37] <= char44_3[37];
                                                  char44_3[38] <= char44_3[38];
                                                  char44_3[39] <= char44_3[39];
                                                  char44_3[40] <= char44_3[40];
                                                  char44_3[41] <= char44_3[41];
                                                  char44_3[42] <= char44_3[42];
                                                  char44_3[43] <= char44_3[43];
                                                  char44_3[44] <= char44_3[44];
                                                  char44_3[45] <= char44_3[45];
                                                  char44_3[46] <= char44_3[46];
                                                  char44_3[47] <= char44_3[47];
                                                  char44_3[48] <= char44_3[48];
                                                  char44_3[49] <= char44_3[49];
                                                  char44_3[50] <= char44_3[50];
                                                  char44_3[51] <= char44_3[51];
                                                  char44_3[52] <= char44_3[52];
                                                  char44_3[53] <= char44_3[53];
                                                  char44_3[54] <= char44_3[54];
                                                  char44_3[55] <= char44_3[55];
                                                  char44_3[56] <= char44_3[56];
                                                  char44_3[57] <= char44_3[57];
                                                  char44_3[58] <= char44_3[58];
                                                  char44_3[59] <= char44_3[59];
                                                  char44_3[60] <= char44_3[60];
                                                  char44_3[61] <= char44_3[61];
                                                  char44_3[62] <= char44_3[62];
                                                  char44_3[63] <= char44_3[63];
                                              end
                                          endcase
                         
                              case((a2 - t1*(a2/t1))/o1)
                                         4'd0: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h000FF000000000000000000000000000;
                                               char44_4[11] <= 128'h003FFC00000000000000000000000000;
                                               char44_4[12] <= 128'h007E7E00800000000000000000000000;
                                               char44_4[13] <= 128'h00F81F00000000000000000000000000;
                                               char44_4[14] <= 128'h01F00F80000000000000000000000000;
                                               char44_4[15] <= 128'h03F00FC0000000000000000000000000;
                                               char44_4[16] <= 128'h03E007C0000000000000000000000000;
                                               char44_4[17] <= 128'h07E007E0000000000000000000000000;
                                               char44_4[18] <= 128'h07C003E0000000000000000000000000;
                                               char44_4[19] <= 128'h0FC003F0000000000000000000000000;
                                               char44_4[20] <= 128'h0FC003F0000000000000000000000000;
                                               char44_4[21] <= 128'h0FC003F0000000000000000000000000;
                                               char44_4[22] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[23] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[24] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[25] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[26] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[27] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[28] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[29] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[30] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[31] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[32] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[33] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[34] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[35] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[36] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[37] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[38] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[39] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[40] <= 128'h1F8001F8000000000000000000000000;
                                               char44_4[41] <= 128'h1F8001F0000000000000000000000000;
                                               char44_4[42] <= 128'h0F8003F0000000000000000000000000;
                                               char44_4[43] <= 128'h0FC003F0000000000000000000000000;
                                               char44_4[44] <= 128'h0FC003F0000000000000000000000000;
                                               char44_4[45] <= 128'h07C003E0000000000000000000000000;
                                               char44_4[46] <= 128'h07E007E0000000000000000000000000;
                                               char44_4[47] <= 128'h03E007C0000000000000000000000000;
                                               char44_4[48] <= 128'h03F00FC0000000000000000000000000;
                                               char44_4[49] <= 128'h01F00F80000000000000000000000000;
                                               char44_4[50] <= 128'h00F81F00000000000000000000000000;
                                               char44_4[51] <= 128'h007E7E00000000000000000000000000;
                                               char44_4[52] <= 128'h003FFC00000000000000000000000000;
                                               char44_4[53] <= 128'h000FF000000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//0
                                         4'd1: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h0000E000000000000000000000000000;
                                               char44_4[11] <= 128'h0001E000000000000000000000000000;
                                               char44_4[12] <= 128'h0003E000000000000000000000000000;
                                               char44_4[13] <= 128'h001FE000000000000000000000000000;
                                               char44_4[14] <= 128'h03FFE000000000000000000000000000;
                                               char44_4[15] <= 128'h03FFE000000000000000000000000000;
                                               char44_4[16] <= 128'h0007E000000000000000000000000000;
                                               char44_4[17] <= 128'h0007E000000000000000000000000000;
                                               char44_4[18] <= 128'h0007E000000000000000000000000000;
                                               char44_4[19] <= 128'h0007E000000000000000000000000000;
                                               char44_4[20] <= 128'h0007E000000000000000000000000000;
                                               char44_4[21] <= 128'h0007E000000000000000000000000000;
                                               char44_4[22] <= 128'h0007E000000000000000000000000000;
                                               char44_4[23] <= 128'h0007E000000000000000000000000000;
                                               char44_4[24] <= 128'h0007E000000000000000000000000000;
                                               char44_4[25] <= 128'h0007E000000000000000000000000000;
                                               char44_4[26] <= 128'h0007E000000000000000000000000000;
                                               char44_4[27] <= 128'h0007E000000000000000000000000000;
                                               char44_4[28] <= 128'h0007E000000000000000000000000000;
                                               char44_4[29] <= 128'h0007E000000000000000000000000000;
                                               char44_4[30] <= 128'h0007E000000000000000000000000000;
                                               char44_4[31] <= 128'h0007E000000000000000000000000000;
                                               char44_4[32] <= 128'h0007E000000000000000000000000000;
                                               char44_4[33] <= 128'h0007E000000000000000000000000000;
                                               char44_4[34] <= 128'h0007E000000000000000000000000000;
                                               char44_4[35] <= 128'h0007E000000000000000000000000000;
                                               char44_4[36] <= 128'h0007E000000000000000000000000000;
                                               char44_4[37] <= 128'h0007E000000000000000000000000000;
                                               char44_4[38] <= 128'h0007E000000000000000000000000000;
                                               char44_4[39] <= 128'h0007E000000000000000000000000000;
                                               char44_4[40] <= 128'h0007E000000000000000000000000000;
                                               char44_4[41] <= 128'h0007E000000000000000000000000000;
                                               char44_4[42] <= 128'h0007E000000000000000000000000000;
                                               char44_4[43] <= 128'h0007E000000000000000000000000000;
                                               char44_4[44] <= 128'h0007E000000000000000000000000000;
                                               char44_4[45] <= 128'h0007E000000000000000000000000000;
                                               char44_4[46] <= 128'h0007E000000000000000000000000000;
                                               char44_4[47] <= 128'h0007E000000000000000000000000000;
                                               char44_4[48] <= 128'h0007E000000000000000000000000000;
                                               char44_4[49] <= 128'h0007E000000000000000000000000000;
                                               char44_4[50] <= 128'h0007E000000000000000000000000000;
                                               char44_4[51] <= 128'h000FF800000000000000000000000000;
                                               char44_4[52] <= 128'h03FFFFC0000000000000000000000000;
                                               char44_4[53] <= 128'h03FFFFC0000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//1
                                         4'd2: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h001FFC00000000000000000000000000;
                                               char44_4[11] <= 128'h007FFF00000000000000000000000000;
                                               char44_4[12] <= 128'h01F83F80000000000000000000000000;
                                               char44_4[13] <= 128'h03E00FC0000000000000000000000000;
                                               char44_4[14] <= 128'h07C007E0000000000000000000000000;
                                               char44_4[15] <= 128'h078007E0000000000000000000000000;
                                               char44_4[16] <= 128'h0F8003F0000000000000000000000000;
                                               char44_4[17] <= 128'h0F8003F0000000000000000000000000;
                                               char44_4[18] <= 128'h1F8003F0000000000000000000000000;
                                               char44_4[19] <= 128'h1F8003F0000000000000000000000000;
                                               char44_4[20] <= 128'h1FC003F0000000000000000000000000;
                                               char44_4[21] <= 128'h1FC003F0000000000000000000000000;
                                               char44_4[22] <= 128'h1FC003F0000000000000000000000000;
                                               char44_4[23] <= 128'h0FC003F0000000000000000000000000;
                                               char44_4[24] <= 128'h07C003F0000000000000000000000000;
                                               char44_4[25] <= 128'h000003E0000000000000000000000000;
                                               char44_4[26] <= 128'h000007E0000000000000000000000000;
                                               char44_4[27] <= 128'h000007E0000000000000000000000000;
                                               char44_4[28] <= 128'h00000FC0000000000000000000000000;
                                               char44_4[29] <= 128'h00000F80000000000000000000000000;
                                               char44_4[30] <= 128'h00001F80000000000000000000000000;
                                               char44_4[31] <= 128'h00003F00000000000000000000000000;
                                               char44_4[32] <= 128'h00003E00000000000000000000000000;
                                               char44_4[33] <= 128'h00007C00000000000000000000000000;
                                               char44_4[34] <= 128'h0000F800000000000000000000000000;
                                               char44_4[35] <= 128'h0001F000000000000000000000000000;
                                               char44_4[36] <= 128'h0003E000000000000000000000000000;
                                               char44_4[37] <= 128'h0007C000000000000000000000000000;
                                               char44_4[38] <= 128'h000F8000000000000000000000000000;
                                               char44_4[39] <= 128'h001F0000000000000000000000000000;
                                               char44_4[40] <= 128'h003E0000000000000000000000000000;
                                               char44_4[41] <= 128'h007C0000000000000000000000000000;
                                               char44_4[42] <= 128'h00F80000000000000000000000000000;
                                               char44_4[43] <= 128'h01F00038000000000000000000000000;
                                               char44_4[44] <= 128'h01E00038000000000000000000000000;
                                               char44_4[45] <= 128'h03C00070000000000000000000000000;
                                               char44_4[46] <= 128'h07800070000000000000000000000000;
                                               char44_4[47] <= 128'h0F8000F0000000000000000000000000;
                                               char44_4[48] <= 128'h0F0000F0000000000000000000000000;
                                               char44_4[49] <= 128'h1E0003F0000000000000000000000000;
                                               char44_4[50] <= 128'h3FFFFFF0000000000000000000000000;
                                               char44_4[51] <= 128'h3FFFFFF0000000000000000000000000;
                                               char44_4[52] <= 128'h3FFFFFE0000000000000000000000000;
                                               char44_4[53] <= 128'h3FFFFFE0000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//2
                                         4'd3: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h003FF000000000000000000000000000;
                                               char44_4[11] <= 128'h00FFFC00000000000000000000000000;
                                               char44_4[12] <= 128'h01F07E00000000000000000000000000;
                                               char44_4[13] <= 128'h03C03F00000000000000000000000000;
                                               char44_4[14] <= 128'h07801F80000000000000000000000000;
                                               char44_4[15] <= 128'h0F800FC0000000000000000000000000;
                                               char44_4[16] <= 128'h0F800FC0000000000000000000000000;
                                               char44_4[17] <= 128'h0F8007E0000000000000000000000000;
                                               char44_4[18] <= 128'h0FC007E0000000000000000000000000;
                                               char44_4[19] <= 128'h0FC007E0000000000000000000000000;
                                               char44_4[20] <= 128'h0FC007E0000000000000000000000000;
                                               char44_4[21] <= 128'h07C007E0000000000000000000000000;
                                               char44_4[22] <= 128'h000007E0000000000000000000000000;
                                               char44_4[23] <= 128'h000007E0000000000000000000000000;
                                               char44_4[24] <= 128'h000007C0000000000000000000000000;
                                               char44_4[25] <= 128'h00000FC0000000000000000000000000;
                                               char44_4[26] <= 128'h00000F80000000000000000000000000;
                                               char44_4[27] <= 128'h00001F00000000000000000000000000;
                                               char44_4[28] <= 128'h00007E00000000000000000000000000;
                                               char44_4[29] <= 128'h0003FC00000000000000000000000000;
                                               char44_4[30] <= 128'h001FF000000000000000000000000000;
                                               char44_4[31] <= 128'h001FFC00000000000000000000000000;
                                               char44_4[32] <= 128'h0000FF00000000000000000000000000;
                                               char44_4[33] <= 128'h00001F80000000000000000000000000;
                                               char44_4[34] <= 128'h00000FC0000000000000000000000000;
                                               char44_4[35] <= 128'h000007E0000000000000000000000000;
                                               char44_4[36] <= 128'h000003E0000000000000000000000000;
                                               char44_4[37] <= 128'h000003F0000000000000000000000000;
                                               char44_4[38] <= 128'h000003F0000000000000000000000000;
                                               char44_4[39] <= 128'h000001F0000000000000000000000000;
                                               char44_4[40] <= 128'h000001F8000000000000000000000000;
                                               char44_4[41] <= 128'h000001F8000000000000000000000000;
                                               char44_4[42] <= 128'h078001F8000000000000000000000000;
                                               char44_4[43] <= 128'h0FC001F8000000000000000000000000;
                                               char44_4[44] <= 128'h1FC001F8000000000000000000000000;
                                               char44_4[45] <= 128'h1FC003F0000000000000000000000000;
                                               char44_4[46] <= 128'h1FC003F0000000000000000000000000;
                                               char44_4[47] <= 128'h1FC003E0000000000000000000000000;
                                               char44_4[48] <= 128'h0F8007E0000000000000000000000000;
                                               char44_4[49] <= 128'h0F8007C0000000000000000000000000;
                                               char44_4[50] <= 128'h07C01F80000000000000000000000000;
                                               char44_4[51] <= 128'h03F07F00000000000000000000000000;
                                               char44_4[52] <= 128'h01FFFE00000000000000000000000000;
                                               char44_4[53] <= 128'h003FF000000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//3
                                         4'd4: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h00001F00000000000000000000000000;
                                               char44_4[11] <= 128'h00001F00000000000000000000000000;
                                               char44_4[12] <= 128'h00003F00000000000000000000000000;
                                               char44_4[13] <= 128'h00003F00000000000000000000000000;
                                               char44_4[14] <= 128'h00007F00000000000000000000000000;
                                               char44_4[15] <= 128'h0000FF00000000000000000000000000;
                                               char44_4[16] <= 128'h0000FF00000000000000000000000000;
                                               char44_4[17] <= 128'h0001FF00000000000000000000000000;
                                               char44_4[18] <= 128'h0003FF00000000000000000000000000;
                                               char44_4[19] <= 128'h0003BF00000000000000000000000000;
                                               char44_4[20] <= 128'h0007BF00000000000000000000000000;
                                               char44_4[21] <= 128'h00073F00000000000000000000000000;
                                               char44_4[22] <= 128'h000F3F00000000000000000000000000;
                                               char44_4[23] <= 128'h001E3F00000000000000000000000000;
                                               char44_4[24] <= 128'h001C3F00000000000000000000000000;
                                               char44_4[25] <= 128'h003C3F00000000000000000000000000;
                                               char44_4[26] <= 128'h00783F00000000000000000000000000;
                                               char44_4[27] <= 128'h00783F00000000000000000000000000;
                                               char44_4[28] <= 128'h00F03F00000000000000000000000000;
                                               char44_4[29] <= 128'h00E03F00000000000000000000000000;
                                               char44_4[30] <= 128'h01E03F00000000000000000000000000;
                                               char44_4[31] <= 128'h03C03F00000000000000000000000000;
                                               char44_4[32] <= 128'h03803F00000000000000000000000000;
                                               char44_4[33] <= 128'h07803F00000000000000000000000000;
                                               char44_4[34] <= 128'h0F003F00000000000000000000000000;
                                               char44_4[35] <= 128'h0F003F00000000000000000000000000;
                                               char44_4[36] <= 128'h1E003F00000000000000000000000000;
                                               char44_4[37] <= 128'h1C003F00000000000000000000000000;
                                               char44_4[38] <= 128'h3C003F00000000000000000000000000;
                                               char44_4[39] <= 128'h7FFFFFFE000000000000000000000000;
                                               char44_4[40] <= 128'h7FFFFFFE000000000000000000000000;
                                               char44_4[41] <= 128'h00003F00000000000000000000000000;
                                               char44_4[42] <= 128'h00003F00000000000000000000000000;
                                               char44_4[43] <= 128'h00003F00000000000000000000000000;
                                               char44_4[44] <= 128'h00003F00000000000000000000000000;
                                               char44_4[45] <= 128'h00003F00000000000000000000000000;
                                               char44_4[46] <= 128'h00003F00000000000000000000000000;
                                               char44_4[47] <= 128'h00003F00000000000000000000000000;
                                               char44_4[48] <= 128'h00003F00000000000000000000000000;
                                               char44_4[49] <= 128'h00003F00000000000000000000000000;
                                               char44_4[50] <= 128'h00003F00000000000000000000000000;
                                               char44_4[51] <= 128'h00007F80000000000000000000000000;
                                               char44_4[52] <= 128'h000FFFFC000000000000000000000000;
                                               char44_4[53] <= 128'h000FFFFC000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//4
                                         4'd5: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h00000000000000000000000000000000;
                                               char44_4[11] <= 128'h03FFFFF0000000000000000000000000;
                                               char44_4[12] <= 128'h03FFFFF0000000000000000000000000;
                                               char44_4[13] <= 128'h03FFFFF0000000000000000000000000;
                                               char44_4[14] <= 128'h03FFFFE0000000000000000000000000;
                                               char44_4[15] <= 128'h03800000000000000000000000000000;
                                               char44_4[16] <= 128'h03800000000000000000000000000000;
                                               char44_4[17] <= 128'h03800000000000000000000000000000;
                                               char44_4[18] <= 128'h03800000000000000000000000000000;
                                               char44_4[19] <= 128'h03800000000000000000000000000000;
                                               char44_4[20] <= 128'h07800000000000000000000000000000;
                                               char44_4[21] <= 128'h07800000000000000000000000000000;
                                               char44_4[22] <= 128'h07800000000000000000000000000000;
                                               char44_4[23] <= 128'h07800000000000000000000000000000;
                                               char44_4[24] <= 128'h07800000000000000000000000000000;
                                               char44_4[25] <= 128'h07800000000000000000000000000000;
                                               char44_4[26] <= 128'h078FF800000000000000000000000000;
                                               char44_4[27] <= 128'h073FFE00000000000000000000000000;
                                               char44_4[28] <= 128'h077FFF80000000000000000000000000;
                                               char44_4[29] <= 128'h07FC3F80000000000000000000000000;
                                               char44_4[30] <= 128'h07E00FC0000000000000000000000000;
                                               char44_4[31] <= 128'h07C007E0000000000000000000000000;
                                               char44_4[32] <= 128'h078007E0000000000000000000000000;
                                               char44_4[33] <= 128'h078003F0000000000000000000000000;
                                               char44_4[34] <= 128'h000003F0000000000000000000000000;
                                               char44_4[35] <= 128'h000001F0000000000000000000000000;
                                               char44_4[36] <= 128'h000001F8000000000000000000000000;
                                               char44_4[37] <= 128'h000001F8000000000000000000000000;
                                               char44_4[38] <= 128'h000001F8000000000000000000000000;
                                               char44_4[39] <= 128'h000001F8000000000000000000000000;
                                               char44_4[40] <= 128'h000001F8000000000000000000000000;
                                               char44_4[41] <= 128'h078001F8000000000000000000000000;
                                               char44_4[42] <= 128'h0FC001F8000000000000000000000000;
                                               char44_4[43] <= 128'h1FC001F0000000000000000000000000;
                                               char44_4[44] <= 128'h1FC001F0000000000000000000000000;
                                               char44_4[45] <= 128'h1FC003F0000000000000000000000000;
                                               char44_4[46] <= 128'h1F8003F0000000000000000000000000;
                                               char44_4[47] <= 128'h1F8003E0000000000000000000000000;
                                               char44_4[48] <= 128'h0F8007E0000000000000000000000000;
                                               char44_4[49] <= 128'h078007C0000000000000000000000000;
                                               char44_4[50] <= 128'h07C01F80000000000000000000000000;
                                               char44_4[51] <= 128'h03F83F00000000000000000000000000;
                                               char44_4[52] <= 128'h00FFFE00000000000000000000000000;
                                               char44_4[53] <= 128'h003FF800000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//5
                                         4'd6: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h0007FE00000000000000000000000000;
                                               char44_4[11] <= 128'h001FFF80000000000000000000000000;
                                               char44_4[12] <= 128'h003F0FC0000000000000000000000000;
                                               char44_4[13] <= 128'h007C07C0000000000000000000000000;
                                               char44_4[14] <= 128'h00F807E0000000000000000000000000;
                                               char44_4[15] <= 128'h01F007E0000000000000000000000000;
                                               char44_4[16] <= 128'h03E007E0000000000000000000000000;
                                               char44_4[17] <= 128'h03C007E0000000000000000000000000;
                                               char44_4[18] <= 128'h07C003C0000000000000000000000000;
                                               char44_4[19] <= 128'h07C00000000000000000000000000000;
                                               char44_4[20] <= 128'h0FC00000000000000000000000000000;
                                               char44_4[21] <= 128'h0F800000000000000000000000000000;
                                               char44_4[22] <= 128'h0F800000000000000000000000000000;
                                               char44_4[23] <= 128'h1F800000000000000000000000000000;
                                               char44_4[24] <= 128'h1F800000000000000000000000000000;
                                               char44_4[25] <= 128'h1F800000000000000000000000000000;
                                               char44_4[26] <= 128'h1F87FE00000000000000000000000000;
                                               char44_4[27] <= 128'h1F9FFF80000000000000000000000000;
                                               char44_4[28] <= 128'h1FBFFFC0000000000000000000000000;
                                               char44_4[29] <= 128'h3FFE1FC0000000000000000000000000;
                                               char44_4[30] <= 128'h3FF807E0000000000000000000000000;
                                               char44_4[31] <= 128'h3FE003F0000000000000000000000000;
                                               char44_4[32] <= 128'h3FE003F0000000000000000000000000;
                                               char44_4[33] <= 128'h3FC001F8000000000000000000000000;
                                               char44_4[34] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[35] <= 128'h3F8001F8000000000000000000000000;
                                               char44_4[36] <= 128'h3F8000F8000000000000000000000000;
                                               char44_4[37] <= 128'h3F8000F8000000000000000000000000;
                                               char44_4[38] <= 128'h3F8000F8000000000000000000000000;
                                               char44_4[39] <= 128'h1F8000F8000000000000000000000000;
                                               char44_4[40] <= 128'h1F8000F8000000000000000000000000;
                                               char44_4[41] <= 128'h1F8000F8000000000000000000000000;
                                               char44_4[42] <= 128'h1F8000F8000000000000000000000000;
                                               char44_4[43] <= 128'h1F8000F8000000000000000000000000;
                                               char44_4[44] <= 128'h0FC001F8000000000000000000000000;
                                               char44_4[45] <= 128'h0FC001F8000000000000000000000000;
                                               char44_4[46] <= 128'h0FC001F0000000000000000000000000;
                                               char44_4[47] <= 128'h07E001F0000000000000000000000000;
                                               char44_4[48] <= 128'h03E003E0000000000000000000000000;
                                               char44_4[49] <= 128'h03F003E0000000000000000000000000;
                                               char44_4[50] <= 128'h01F807C0000000000000000000000000;
                                               char44_4[51] <= 128'h00FE1F80000000000000000000000000;
                                               char44_4[52] <= 128'h007FFE00000000000000000000000000;
                                               char44_4[53] <= 128'h001FF800000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//6
                                         4'd7: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h00000000000000000000000000000000;
                                               char44_4[11] <= 128'h07FFFFF8000000000000000000000000;
                                               char44_4[12] <= 128'h07FFFFF8000000000000000000000000;
                                               char44_4[13] <= 128'h07FFFFF8000000000000000000000000;
                                               char44_4[14] <= 128'h0FFFFFF0000000000000000000000000;
                                               char44_4[15] <= 128'h0FC000E0000000000000000000000000;
                                               char44_4[16] <= 128'h0F8001E0000000000000000000000000;
                                               char44_4[17] <= 128'h0F0001C0000000000000000000000000;
                                               char44_4[18] <= 128'h0E0003C0000000000000000000000000;
                                               char44_4[19] <= 128'h0E000780000000000000000000000000;
                                               char44_4[20] <= 128'h1E000780000000000000000000000000;
                                               char44_4[21] <= 128'h1C000F00000000000000000000000000;
                                               char44_4[22] <= 128'h00000F00000000000000000000000000;
                                               char44_4[23] <= 128'h00001E00000000000000000000000000;
                                               char44_4[24] <= 128'h00001E00000000000000000000000000;
                                               char44_4[25] <= 128'h00003C00000000000000000000000000;
                                               char44_4[26] <= 128'h00003C00000000000000000000000000;
                                               char44_4[27] <= 128'h00007800000000000000000000000000;
                                               char44_4[28] <= 128'h00007800000000000000000000000000;
                                               char44_4[29] <= 128'h0000F800000000000000000000000000;
                                               char44_4[30] <= 128'h0000F000000000000000000000000000;
                                               char44_4[31] <= 128'h0001F000000000000000000000000000;
                                               char44_4[32] <= 128'h0001E000000000000000000000000000;
                                               char44_4[33] <= 128'h0003E000000000000000000000000000;
                                               char44_4[34] <= 128'h0003E000000000000000000000000000;
                                               char44_4[35] <= 128'h0003E000000000000000000000000000;
                                               char44_4[36] <= 128'h0007C000000000000000000000000000;
                                               char44_4[37] <= 128'h0007C000000000000000000000000000;
                                               char44_4[38] <= 128'h0007C000000000000000000000000000;
                                               char44_4[39] <= 128'h000FC000000000000000000000000000;
                                               char44_4[40] <= 128'h000FC000000000000000000000000000;
                                               char44_4[41] <= 128'h000FC000000000000000000000000000;
                                               char44_4[42] <= 128'h000FC000000000000000000000000000;
                                               char44_4[43] <= 128'h001FC000000000000000000000000000;
                                               char44_4[44] <= 128'h001FC000000000000000000000000000;
                                               char44_4[45] <= 128'h001FC000000000000000000000000000;
                                               char44_4[46] <= 128'h001FC000000000000000000000000000;
                                               char44_4[47] <= 128'h001FC000000000000000000000000000;
                                               char44_4[48] <= 128'h001FC000000000000000000000000000;
                                               char44_4[49] <= 128'h001FC000000000000000000000000000;
                                               char44_4[50] <= 128'h001FC000000000000000000000000000;
                                               char44_4[51] <= 128'h001FC000000000000000000000000000;
                                               char44_4[52] <= 128'h001FC000000000000000000000000000;
                                               char44_4[53] <= 128'h000F8000000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//7
                                         4'd8: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h003FF800000000000000000000000000;
                                               char44_4[11] <= 128'h00FFFE00000000000000000000000000;
                                               char44_4[12] <= 128'h01F81F80000000000000000000000000;
                                               char44_4[13] <= 128'h03E00FC0000000000000000000000000;
                                               char44_4[14] <= 128'h07C003E0000000000000000000000000;
                                               char44_4[15] <= 128'h0F8003E0000000000000000000000000;
                                               char44_4[16] <= 128'h0F8001F0000000000000000000000000;
                                               char44_4[17] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[18] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[19] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[20] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[21] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[22] <= 128'h1F8001F0000000000000000000000000;
                                               char44_4[23] <= 128'h1FC001F0000000000000000000000000;
                                               char44_4[24] <= 128'h0FC001F0000000000000000000000000;
                                               char44_4[25] <= 128'h0FF003E0000000000000000000000000;
                                               char44_4[26] <= 128'h07F803C0000000000000000000000000;
                                               char44_4[27] <= 128'h03FE0F80000000000000000000000000;
                                               char44_4[28] <= 128'h01FF9F00000000000000000000000000;
                                               char44_4[29] <= 128'h00FFFE00000000000000000000000000;
                                               char44_4[30] <= 128'h003FF800000000000000000000000000;
                                               char44_4[31] <= 128'h007FFC00000000000000000000000000;
                                               char44_4[32] <= 128'h01F7FF00000000000000000000000000;
                                               char44_4[33] <= 128'h03E1FF80000000000000000000000000;
                                               char44_4[34] <= 128'h07C07FC0000000000000000000000000;
                                               char44_4[35] <= 128'h0F801FE0000000000000000000000000;
                                               char44_4[36] <= 128'h0F800FE0000000000000000000000000;
                                               char44_4[37] <= 128'h1F0007F0000000000000000000000000;
                                               char44_4[38] <= 128'h1F0003F0000000000000000000000000;
                                               char44_4[39] <= 128'h3E0001F8000000000000000000000000;
                                               char44_4[40] <= 128'h3E0001F8000000000000000000000000;
                                               char44_4[41] <= 128'h3E0001F8000000000000000000000000;
                                               char44_4[42] <= 128'h3E0000F8000000000000000000000000;
                                               char44_4[43] <= 128'h3E0000F8000000000000000000000000;
                                               char44_4[44] <= 128'h3E0000F8000000000000000000000000;
                                               char44_4[45] <= 128'h3E0000F8000000000000000000000000;
                                               char44_4[46] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[47] <= 128'h1F0001F0000000000000000000000000;
                                               char44_4[48] <= 128'h0F8003E0000000000000000000000000;
                                               char44_4[49] <= 128'h0FC003E0000000000000000000000000;
                                               char44_4[50] <= 128'h07E007C0000000000000000000000000;
                                               char44_4[51] <= 128'h01F83F80000000000000000000000000;
                                               char44_4[52] <= 128'h00FFFE00000000000000000000000000;
                                               char44_4[53] <= 128'h003FF800000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//8
                                         4'd9: begin
                                               char44_4[0] <= 128'h00000000000000000000000000000000;
                                               char44_4[1] <= 128'h00000000000000000000000000000000;
                                               char44_4[2] <= 128'h00000000000000000000000000000000;
                                               char44_4[3] <= 128'h00000000000000000000000000000000;
                                               char44_4[4] <= 128'h00000000000000000000000000000000;
                                               char44_4[5] <= 128'h00000000000000000000000000000000;
                                               char44_4[6] <= 128'h00000000000000000000000000000000;
                                               char44_4[7] <= 128'h00000000000000000000000000000000;
                                               char44_4[8] <= 128'h00000000000000000000000000000000;
                                               char44_4[9] <= 128'h00000000000000000000000000000000;
                                               char44_4[10] <= 128'h003FF000000000000000000000000000;
                                               char44_4[11] <= 128'h00FFFC00000000000000000000000000;
                                               char44_4[12] <= 128'h01F83F00000000000000000000000000;
                                               char44_4[13] <= 128'h03E01F80000000000000000000000000;
                                               char44_4[14] <= 128'h07C00F80000000000000000000000000;
                                               char44_4[15] <= 128'h0FC007C0000000000000000000000000;
                                               char44_4[16] <= 128'h0F8003E0000000000000000000000000;
                                               char44_4[17] <= 128'h1F8003E0000000000000000000000000;
                                               char44_4[18] <= 128'h1F0003F0000000000000000000000000;
                                               char44_4[19] <= 128'h1F0003F0000000000000000000000000;
                                               char44_4[20] <= 128'h3F0001F0000000000000000000000000;
                                               char44_4[21] <= 128'h3F0001F0000000000000000000000000;
                                               char44_4[22] <= 128'h3F0001F8000000000000000000000000;
                                               char44_4[23] <= 128'h3F0001F8000000000000000000000000;
                                               char44_4[24] <= 128'h3F0001F8000000000000000000000000;
                                               char44_4[25] <= 128'h3F0001F8000000000000000000000000;
                                               char44_4[26] <= 128'h3F0001F8000000000000000000000000;
                                               char44_4[27] <= 128'h3F0001F8000000000000000000000000;
                                               char44_4[28] <= 128'h3F0003F8000000000000000000000000;
                                               char44_4[29] <= 128'h1F8003F8000000000000000000000000;
                                               char44_4[30] <= 128'h1F8007F8000000000000000000000000;
                                               char44_4[31] <= 128'h1F800FF8000000000000000000000000;
                                               char44_4[32] <= 128'h0FC01FF8000000000000000000000000;
                                               char44_4[33] <= 128'h0FE03FF8000000000000000000000000;
                                               char44_4[34] <= 128'h07F8FDF8000000000000000000000000;
                                               char44_4[35] <= 128'h03FFF9F8000000000000000000000000;
                                               char44_4[36] <= 128'h01FFF1F8000000000000000000000000;
                                               char44_4[37] <= 128'h003F83F8000000000000000000000000;
                                               char44_4[38] <= 128'h000003F0000000000000000000000000;
                                               char44_4[39] <= 128'h000003F0000000000000000000000000;
                                               char44_4[40] <= 128'h000003F0000000000000000000000000;
                                               char44_4[41] <= 128'h000003F0000000000000000000000000;
                                               char44_4[42] <= 128'h000007E0000000000000000000000000;
                                               char44_4[43] <= 128'h000007E0000000000000000000000000;
                                               char44_4[44] <= 128'h000007C0000000000000000000000000;
                                               char44_4[45] <= 128'h03C007C0000000000000000000000000;
                                               char44_4[46] <= 128'h07C00F80000000000000000000000000;
                                               char44_4[47] <= 128'h0FE00F80000000000000000000000000;
                                               char44_4[48] <= 128'h0FE01F00000000000000000000000000;
                                               char44_4[49] <= 128'h0FE03E00000000000000000000000000;
                                               char44_4[50] <= 128'h07E07E00000000000000000000000000;
                                               char44_4[51] <= 128'h07F1F800000000000000000000000000;
                                               char44_4[52] <= 128'h03FFF000000000000000000000000000;
                                               char44_4[53] <= 128'h00FFC000000000000000000000000000;
                                               char44_4[54] <= 128'h00000000000000000000000000000000;
                                               char44_4[55] <= 128'h00000000000000000000000000000000;
                                               char44_4[56] <= 128'h00000000000000000000000000000000;
                                               char44_4[57] <= 128'h00000000000000000000000000000000;
                                               char44_4[58] <= 128'h00000000000000000000000000000000;
                                               char44_4[59] <= 128'h00000000000000000000000000000000;
                                               char44_4[60] <= 128'h00000000000000000000000000000000;
                                               char44_4[61] <= 128'h00000000000000000000000000000000;
                                               char44_4[62] <= 128'h00000000000000000000000000000000;
                                               char44_4[63] <= 128'h00000000000000000000000000000000;
                                         end//9
                                         default: begin
                                             char44_4[0] <= char44_4[0];
                                             char44_4[1] <= char44_4[1];
                                             char44_4[2] <= char44_4[2];
                                             char44_4[3] <= char44_4[3];
                                             char44_4[4] <= char44_4[4];
                                             char44_4[5] <= char44_4[5];
                                             char44_4[6] <= char44_4[6];
                                             char44_4[7] <= char44_4[7];
                                             char44_4[8] <= char44_4[8];
                                             char44_4[9] <= char44_4[9];
                                             char44_4[10] <= char44_4[10];
                                             char44_4[11] <= char44_4[11];
                                             char44_4[12] <= char44_4[12];
                                             char44_4[13] <= char44_4[13];
                                             char44_4[14] <= char44_4[14];
                                             char44_4[15] <= char44_4[15];
                                             char44_4[16] <= char44_4[16];
                                             char44_4[17] <= char44_4[17];
                                             char44_4[18] <= char44_4[18];
                                             char44_4[19] <= char44_4[19];
                                             char44_4[20] <= char44_4[20];
                                             char44_4[21] <= char44_4[21];
                                             char44_4[22] <= char44_4[22];
                                             char44_4[23] <= char44_4[23];
                                             char44_4[24] <= char44_4[24];
                                             char44_4[25] <= char44_4[25];
                                             char44_4[26] <= char44_4[26];
                                             char44_4[27] <= char44_4[27];
                                             char44_4[28] <= char44_4[28];
                                             char44_4[29] <= char44_4[29];
                                             char44_4[30] <= char44_4[30];
                                             char44_4[31] <= char44_4[31];
                                             char44_4[32] <= char44_4[32];
                                             char44_4[33] <= char44_4[33];
                                             char44_4[34] <= char44_4[34];
                                             char44_4[35] <= char44_4[35];
                                             char44_4[36] <= char44_4[36];
                                             char44_4[37] <= char44_4[37];
                                             char44_4[38] <= char44_4[38];
                                             char44_4[39] <= char44_4[39];
                                             char44_4[40] <= char44_4[40];
                                             char44_4[41] <= char44_4[41];
                                             char44_4[42] <= char44_4[42];
                                             char44_4[43] <= char44_4[43];
                                             char44_4[44] <= char44_4[44];
                                             char44_4[45] <= char44_4[45];
                                             char44_4[46] <= char44_4[46];
                                             char44_4[47] <= char44_4[47];
                                             char44_4[48] <= char44_4[48];
                                             char44_4[49] <= char44_4[49];
                                             char44_4[50] <= char44_4[50];
                                             char44_4[51] <= char44_4[51];
                                             char44_4[52] <= char44_4[52];
                                             char44_4[53] <= char44_4[53];
                                             char44_4[54] <= char44_4[54];
                                             char44_4[55] <= char44_4[55];
                                             char44_4[56] <= char44_4[56];
                                             char44_4[57] <= char44_4[57];
                                             char44_4[58] <= char44_4[58];
                                             char44_4[59] <= char44_4[59];
                                             char44_4[60] <= char44_4[60];
                                             char44_4[61] <= char44_4[61];
                                             char44_4[62] <= char44_4[62];
                                             char44_4[63] <= char44_4[63];
                                         end
                                     endcase
                             

    char[  0] <= {char22_0[0], char22_1[0], char22_2[0], char22_3[0], char22_4[0], char2[0]};
    char[  1] <= {char22_0[1], char22_1[1], char22_2[1], char22_3[1], char22_4[1], char2[1]};
    char[  2] <= {char22_0[2], char22_1[2], char22_2[2], char22_3[2], char22_4[2], char2[2]};
    char[  3] <= {char22_0[3], char22_1[3], char22_2[3], char22_3[3], char22_4[3], char2[3]};
    char[  4] <= {char22_0[4], char22_1[4], char22_2[4], char22_3[4], char22_4[4], char2[4]};
    char[  5] <= {char22_0[5], char22_1[5], char22_2[5], char22_3[5], char22_4[5], char2[5]};
    char[  6] <= {char22_0[6], char22_1[6], char22_2[6], char22_3[6], char22_4[6], char2[6]};
    char[  7] <= {char22_0[7], char22_1[7], char22_2[7], char22_3[7], char22_4[7], char2[7]};
    char[  8] <= {char22_0[8], char22_1[8], char22_2[8], char22_3[8], char22_4[8], char2[8]};
    char[  9] <= {char22_0[9], char22_1[9], char22_2[9], char22_3[9], char22_4[9], char2[9]};
    char[ 10] <= {char22_0[10], char22_1[10], char22_2[10], char22_3[10], char22_4[10], char2[10]};
    char[ 11] <= {char22_0[11], char22_1[11], char22_2[11], char22_3[11], char22_4[11], char2[11]};
    char[ 12] <= {char22_0[12], char22_1[12], char22_2[12], char22_3[12], char22_4[12], char2[12]};
    char[ 13] <= {char22_0[13], char22_1[13], char22_2[13], char22_3[13], char22_4[13], char2[13]};
    char[ 14] <= {char22_0[14], char22_1[14], char22_2[14], char22_3[14], char22_4[14], char2[14]};
    char[ 15] <= {char22_0[15], char22_1[15], char22_2[15], char22_3[15], char22_4[15], char2[15]};
    char[ 16] <= {char22_0[16], char22_1[16], char22_2[16], char22_3[16], char22_4[16], char2[16]};
    char[ 17] <= {char22_0[17], char22_1[17], char22_2[17], char22_3[17], char22_4[17], char2[17]};
    char[ 18] <= {char22_0[18], char22_1[18], char22_2[18], char22_3[18], char22_4[18], char2[18]};
    char[ 19] <= {char22_0[19], char22_1[19], char22_2[19], char22_3[19], char22_4[19], char2[19]};
    char[ 20] <= {char22_0[20], char22_1[20], char22_2[20], char22_3[20], char22_4[20], char2[20]};
    char[ 21] <= {char22_0[21], char22_1[21], char22_2[21], char22_3[21], char22_4[21], char2[21]};
    char[ 22] <= {char22_0[22], char22_1[22], char22_2[22], char22_3[22], char22_4[22], char2[22]};
    char[ 23] <= {char22_0[23], char22_1[23], char22_2[23], char22_3[23], char22_4[23], char2[23]};
    char[ 24] <= {char22_0[24], char22_1[24], char22_2[24], char22_3[24], char22_4[24], char2[24]};
    char[ 25] <= {char22_0[25], char22_1[25], char22_2[25], char22_3[25], char22_4[25], char2[25]};
    char[ 26] <= {char22_0[26], char22_1[26], char22_2[26], char22_3[26], char22_4[26], char2[26]};
    char[ 27] <= {char22_0[27], char22_1[27], char22_2[27], char22_3[27], char22_4[27], char2[27]};
    char[ 28] <= {char22_0[28], char22_1[28], char22_2[28], char22_3[28], char22_4[28], char2[28]};
    char[ 29] <= {char22_0[29], char22_1[29], char22_2[29], char22_3[29], char22_4[29], char2[29]};
    char[ 30] <= {char22_0[30], char22_1[30], char22_2[30], char22_3[30], char22_4[30], char2[30]};
    char[ 31] <= {char22_0[31], char22_1[31], char22_2[31], char22_3[31], char22_4[31], char2[31]};
    char[ 32] <= {char22_0[32], char22_1[32], char22_2[32], char22_3[32], char22_4[32], char2[32]};
    char[ 33] <= {char22_0[33], char22_1[33], char22_2[33], char22_3[33], char22_4[33], char2[33]};
    char[ 34] <= {char22_0[34], char22_1[34], char22_2[34], char22_3[34], char22_4[34], char2[34]};
    char[ 35] <= {char22_0[35], char22_1[35], char22_2[35], char22_3[35], char22_4[35], char2[35]};
    char[ 36] <= {char22_0[36], char22_1[36], char22_2[36], char22_3[36], char22_4[36], char2[36]};
    char[ 37] <= {char22_0[37], char22_1[37], char22_2[37], char22_3[37], char22_4[37], char2[37]};
    char[ 38] <= {char22_0[38], char22_1[38], char22_2[38], char22_3[38], char22_4[38], char2[38]};
    char[ 39] <= {char22_0[39], char22_1[39], char22_2[39], char22_3[39], char22_4[39], char2[39]};
    char[ 40] <= {char22_0[40], char22_1[40], char22_2[40], char22_3[40], char22_4[40], char2[40]};
    char[ 41] <= {char22_0[41], char22_1[41], char22_2[41], char22_3[41], char22_4[41], char2[41]};
    char[ 42] <= {char22_0[42], char22_1[42], char22_2[42], char22_3[42], char22_4[42], char2[42]};
    char[ 43] <= {char22_0[43], char22_1[43], char22_2[43], char22_3[43], char22_4[43], char2[43]};
    char[ 44] <= {char22_0[44], char22_1[44], char22_2[44], char22_3[44], char22_4[44], char2[44]};
    char[ 45] <= {char22_0[45], char22_1[45], char22_2[45], char22_3[45], char22_4[45], char2[45]};
    char[ 46] <= {char22_0[46], char22_1[46], char22_2[46], char22_3[46], char22_4[46], char2[46]};
    char[ 47] <= {char22_0[47], char22_1[47], char22_2[47], char22_3[47], char22_4[47], char2[47]};
    char[ 48] <= {char22_0[48], char22_1[48], char22_2[48], char22_3[48], char22_4[48], char2[48]};
    char[ 49] <= {char22_0[49], char22_1[49], char22_2[49], char22_3[49], char22_4[49], char2[49]};
    char[ 50] <= {char22_0[50], char22_1[50], char22_2[50], char22_3[50], char22_4[50], char2[50]};
    char[ 51] <= {char22_0[51], char22_1[51], char22_2[51], char22_3[51], char22_4[51], char2[51]};
    char[ 52] <= {char22_0[52], char22_1[52], char22_2[52], char22_3[52], char22_4[52], char2[52]};
    char[ 53] <= {char22_0[53], char22_1[53], char22_2[53], char22_3[53], char22_4[53], char2[53]};
    char[ 54] <= {char22_0[54], char22_1[54], char22_2[54], char22_3[54], char22_4[54], char2[54]};
    char[ 55] <= {char22_0[55], char22_1[55], char22_2[55], char22_3[55], char22_4[55], char2[55]};
    char[ 56] <= {char22_0[56], char22_1[56], char22_2[56], char22_3[56], char22_4[56], char2[56]};
    char[ 57] <= {char22_0[57], char22_1[57], char22_2[57], char22_3[57], char22_4[57], char2[57]};
    char[ 58] <= {char22_0[58], char22_1[58], char22_2[58], char22_3[58], char22_4[58], char2[58]};
    char[ 59] <= {char22_0[59], char22_1[59], char22_2[59], char22_3[59], char22_4[59], char2[59]};
    char[ 60] <= {char22_0[60], char22_1[60], char22_2[60], char22_3[60], char22_4[60], char2[60]};
    char[ 61] <= {char22_0[61], char22_1[61], char22_2[61], char22_3[61], char22_4[61], char2[61]};
    char[ 62] <= {char22_0[62], char22_1[62], char22_2[62], char22_3[62], char22_4[62], char2[62]};
    char[ 63] <= {char22_0[63], char22_1[63], char22_2[63], char22_3[63], char22_4[63], char2[63]};
    char[ 64] <= {char33_0[0], char33_1[0], char33_2[0], char33_3[0], char33_4[0], char3[0]};
    char[ 65] <= {char33_0[1], char33_1[1], char33_2[1], char33_3[1], char33_4[1], char3[1]};
    char[ 66] <= {char33_0[2], char33_1[2], char33_2[2], char33_3[2], char33_4[2], char3[2]};
    char[ 67] <= {char33_0[3], char33_1[3], char33_2[3], char33_3[3], char33_4[3], char3[3]};
    char[ 68] <= {char33_0[4], char33_1[4], char33_2[4], char33_3[4], char33_4[4], char3[4]};
    char[ 69] <= {char33_0[5], char33_1[5], char33_2[5], char33_3[5], char33_4[5], char3[5]};
    char[ 70] <= {char33_0[6], char33_1[6], char33_2[6], char33_3[6], char33_4[6], char3[6]};
    char[ 71] <= {char33_0[7], char33_1[7], char33_2[7], char33_3[7], char33_4[7], char3[7]};
    char[ 72] <= {char33_0[8], char33_1[8], char33_2[8], char33_3[8], char33_4[8], char3[8]};
    char[ 73] <= {char33_0[9], char33_1[9], char33_2[9], char33_3[9], char33_4[9], char3[9]};
    char[ 74] <= {char33_0[10], char33_1[10], char33_2[10], char33_3[10], char33_4[10], char3[10]};
    char[ 75] <= {char33_0[11], char33_1[11], char33_2[11], char33_3[11], char33_4[11], char3[11]};
    char[ 76] <= {char33_0[12], char33_1[12], char33_2[12], char33_3[12], char33_4[12], char3[12]};
    char[ 77] <= {char33_0[13], char33_1[13], char33_2[13], char33_3[13], char33_4[13], char3[13]};
    char[ 78] <= {char33_0[14], char33_1[14], char33_2[14], char33_3[14], char33_4[14], char3[14]};
    char[ 79] <= {char33_0[15], char33_1[15], char33_2[15], char33_3[15], char33_4[15], char3[15]};
    char[ 80] <= {char33_0[16], char33_1[16], char33_2[16], char33_3[16], char33_4[16], char3[16]};
    char[ 81] <= {char33_0[17], char33_1[17], char33_2[17], char33_3[17], char33_4[17], char3[17]};
    char[ 82] <= {char33_0[18], char33_1[18], char33_2[18], char33_3[18], char33_4[18], char3[18]};
    char[ 83] <= {char33_0[19], char33_1[19], char33_2[19], char33_3[19], char33_4[19], char3[19]};
    char[ 84] <= {char33_0[20], char33_1[20], char33_2[20], char33_3[20], char33_4[20], char3[20]};
    char[ 85] <= {char33_0[21], char33_1[21], char33_2[21], char33_3[21], char33_4[21], char3[21]};
    char[ 86] <= {char33_0[22], char33_1[22], char33_2[22], char33_3[22], char33_4[22], char3[22]};
    char[ 87] <= {char33_0[23], char33_1[23], char33_2[23], char33_3[23], char33_4[23], char3[23]};
    char[ 88] <= {char33_0[24], char33_1[24], char33_2[24], char33_3[24], char33_4[24], char3[24]};
    char[ 89] <= {char33_0[25], char33_1[25], char33_2[25], char33_3[25], char33_4[25], char3[25]};
    char[ 90] <= {char33_0[26], char33_1[26], char33_2[26], char33_3[26], char33_4[26], char3[26]};
    char[ 91] <= {char33_0[27], char33_1[27], char33_2[27], char33_3[27], char33_4[27], char3[27]};
    char[ 92] <= {char33_0[28], char33_1[28], char33_2[28], char33_3[28], char33_4[28], char3[28]};
    char[ 93] <= {char33_0[29], char33_1[29], char33_2[29], char33_3[29], char33_4[29], char3[29]};
    char[ 94] <= {char33_0[30], char33_1[30], char33_2[30], char33_3[30], char33_4[30], char3[30]};
    char[ 95] <= {char33_0[31], char33_1[31], char33_2[31], char33_3[31], char33_4[31], char3[31]};
    char[ 96] <= {char33_0[32], char33_1[32], char33_2[32], char33_3[32], char33_4[32], char3[32]};
    char[ 97] <= {char33_0[33], char33_1[33], char33_2[33], char33_3[33], char33_4[33], char3[33]};
    char[ 98] <= {char33_0[34], char33_1[34], char33_2[34], char33_3[34], char33_4[34], char3[34]};
    char[ 99] <= {char33_0[35], char33_1[35], char33_2[35], char33_3[35], char33_4[35], char3[35]};
    char[100] <= {char33_0[36], char33_1[36], char33_2[36], char33_3[36], char33_4[36], char3[36]};
    char[101] <= {char33_0[37], char33_1[37], char33_2[37], char33_3[37], char33_4[37], char3[37]};
    char[102] <= {char33_0[38], char33_1[38], char33_2[38], char33_3[38], char33_4[38], char3[38]};
    char[103] <= {char33_0[39], char33_1[39], char33_2[39], char33_3[39], char33_4[39], char3[39]};
    char[104] <= {char33_0[40], char33_1[40], char33_2[40], char33_3[40], char33_4[40], char3[40]};
    char[105] <= {char33_0[41], char33_1[41], char33_2[41], char33_3[41], char33_4[41], char3[41]};
    char[106] <= {char33_0[42], char33_1[42], char33_2[42], char33_3[42], char33_4[42], char3[42]};
    char[107] <= {char33_0[43], char33_1[43], char33_2[43], char33_3[43], char33_4[43], char3[43]};
    char[108] <= {char33_0[44], char33_1[44], char33_2[44], char33_3[44], char33_4[44], char3[44]};
    char[109] <= {char33_0[45], char33_1[45], char33_2[45], char33_3[45], char33_4[45], char3[45]};
    char[110] <= {char33_0[46], char33_1[46], char33_2[46], char33_3[46], char33_4[46], char3[46]};
    char[111] <= {char33_0[47], char33_1[47], char33_2[47], char33_3[47], char33_4[47], char3[47]};
    char[112] <= {char33_0[48], char33_1[48], char33_2[48], char33_3[48], char33_4[48], char3[48]};
    char[113] <= {char33_0[49], char33_1[49], char33_2[49], char33_3[49], char33_4[49], char3[49]};
    char[114] <= {char33_0[50], char33_1[50], char33_2[50], char33_3[50], char33_4[50], char3[50]};
    char[115] <= {char33_0[51], char33_1[51], char33_2[51], char33_3[51], char33_4[51], char3[51]};
    char[116] <= {char33_0[52], char33_1[52], char33_2[52], char33_3[52], char33_4[52], char3[52]};
    char[117] <= {char33_0[53], char33_1[53], char33_2[53], char33_3[53], char33_4[53], char3[53]};
    char[118] <= {char33_0[54], char33_1[54], char33_2[54], char33_3[54], char33_4[54], char3[54]};
    char[119] <= {char33_0[55], char33_1[55], char33_2[55], char33_3[55], char33_4[55], char3[55]};
    char[120] <= {char33_0[56], char33_1[56], char33_2[56], char33_3[56], char33_4[56], char3[56]};
    char[121] <= {char33_0[57], char33_1[57], char33_2[57], char33_3[57], char33_4[57], char3[57]};
    char[122] <= {char33_0[58], char33_1[58], char33_2[58], char33_3[58], char33_4[58], char3[58]};
    char[123] <= {char33_0[59], char33_1[59], char33_2[59], char33_3[59], char33_4[59], char3[59]};
    char[124] <= {char33_0[60], char33_1[60], char33_2[60], char33_3[60], char33_4[60], char3[60]};
    char[125] <= {char33_0[61], char33_1[61], char33_2[61], char33_3[61], char33_4[61], char3[61]};
    char[126] <= {char33_0[62], char33_1[62], char33_2[62], char33_3[62], char33_4[62], char3[62]};
    char[127] <= {char33_0[63], char33_1[63], char33_2[63], char33_3[63], char33_4[63], char3[63]};
    char[128] <= {char44_0[0], char44_1[0], char44_2[0], char44_3[0], char44_4[0], char4[0]};
    char[129] <= {char44_0[1], char44_1[1], char44_2[1], char44_3[1], char44_4[1], char4[1]};
    char[130] <= {char44_0[2], char44_1[2], char44_2[2], char44_3[2], char44_4[2], char4[2]};
    char[131] <= {char44_0[3], char44_1[3], char44_2[3], char44_3[3], char44_4[3], char4[3]};
    char[132] <= {char44_0[4], char44_1[4], char44_2[4], char44_3[4], char44_4[4], char4[4]};
    char[133] <= {char44_0[5], char44_1[5], char44_2[5], char44_3[5], char44_4[5], char4[5]};
    char[134] <= {char44_0[6], char44_1[6], char44_2[6], char44_3[6], char44_4[6], char4[6]};
    char[135] <= {char44_0[7], char44_1[7], char44_2[7], char44_3[7], char44_4[7], char4[7]};
    char[136] <= {char44_0[8], char44_1[8], char44_2[8], char44_3[8], char44_4[8], char4[8]};
    char[137] <= {char44_0[9], char44_1[9], char44_2[9], char44_3[9], char44_4[9], char4[9]};
    char[138] <= {char44_0[10], char44_1[10], char44_2[10], char44_3[10], char44_4[10], char4[10]};
    char[139] <= {char44_0[11], char44_1[11], char44_2[11], char44_3[11], char44_4[11], char4[11]};
    char[140] <= {char44_0[12], char44_1[12], char44_2[12], char44_3[12], char44_4[12], char4[12]};
    char[141] <= {char44_0[13], char44_1[13], char44_2[13], char44_3[13], char44_4[13], char4[13]};
    char[142] <= {char44_0[14], char44_1[14], char44_2[14], char44_3[14], char44_4[14], char4[14]};
    char[143] <= {char44_0[15], char44_1[15], char44_2[15], char44_3[15], char44_4[15], char4[15]};
    char[144] <= {char44_0[16], char44_1[16], char44_2[16], char44_3[16], char44_4[16], char4[16]};
    char[145] <= {char44_0[17], char44_1[17], char44_2[17], char44_3[17], char44_4[17], char4[17]};
    char[146] <= {char44_0[18], char44_1[18], char44_2[18], char44_3[18], char44_4[18], char4[18]};
    char[147] <= {char44_0[19], char44_1[19], char44_2[19], char44_3[19], char44_4[19], char4[19]};
    char[148] <= {char44_0[20], char44_1[20], char44_2[20], char44_3[20], char44_4[20], char4[20]};
    char[149] <= {char44_0[21], char44_1[21], char44_2[21], char44_3[21], char44_4[21], char4[21]};
    char[150] <= {char44_0[22], char44_1[22], char44_2[22], char44_3[22], char44_4[22], char4[22]};
    char[151] <= {char44_0[23], char44_1[23], char44_2[23], char44_3[23], char44_4[23], char4[23]};
    char[152] <= {char44_0[24], char44_1[24], char44_2[24], char44_3[24], char44_4[24], char4[24]};
    char[153] <= {char44_0[25], char44_1[25], char44_2[25], char44_3[25], char44_4[25], char4[25]};
    char[154] <= {char44_0[26], char44_1[26], char44_2[26], char44_3[26], char44_4[26], char4[26]};
    char[155] <= {char44_0[27], char44_1[27], char44_2[27], char44_3[27], char44_4[27], char4[27]};
    char[156] <= {char44_0[28], char44_1[28], char44_2[28], char44_3[28], char44_4[28], char4[28]};
    char[157] <= {char44_0[29], char44_1[29], char44_2[29], char44_3[29], char44_4[29], char4[29]};
    char[158] <= {char44_0[30], char44_1[30], char44_2[30], char44_3[30], char44_4[30], char4[30]};
    char[159] <= {char44_0[31], char44_1[31], char44_2[31], char44_3[31], char44_4[31], char4[31]};
    char[160] <= {char44_0[32], char44_1[32], char44_2[32], char44_3[32], char44_4[32], char4[32]};
    char[161] <= {char44_0[33], char44_1[33], char44_2[33], char44_3[33], char44_4[33], char4[33]};
    char[162] <= {char44_0[34], char44_1[34], char44_2[34], char44_3[34], char44_4[34], char4[34]};
    char[163] <= {char44_0[35], char44_1[35], char44_2[35], char44_3[35], char44_4[35], char4[35]};
    char[164] <= {char44_0[36], char44_1[36], char44_2[36], char44_3[36], char44_4[36], char4[36]};
    char[165] <= {char44_0[37], char44_1[37], char44_2[37], char44_3[37], char44_4[37], char4[37]};
    char[166] <= {char44_0[38], char44_1[38], char44_2[38], char44_3[38], char44_4[38], char4[38]};
    char[167] <= {char44_0[39], char44_1[39], char44_2[39], char44_3[39], char44_4[39], char4[39]};
    char[168] <= {char44_0[40], char44_1[40], char44_2[40], char44_3[40], char44_4[40], char4[40]};
    char[169] <= {char44_0[41], char44_1[41], char44_2[41], char44_3[41], char44_4[41], char4[41]};
    char[170] <= {char44_0[42], char44_1[42], char44_2[42], char44_3[42], char44_4[42], char4[42]};
    char[171] <= {char44_0[43], char44_1[43], char44_2[43], char44_3[43], char44_4[43], char4[43]};
    char[172] <= {char44_0[44], char44_1[44], char44_2[44], char44_3[44], char44_4[44], char4[44]};
    char[173] <= {char44_0[45], char44_1[45], char44_2[45], char44_3[45], char44_4[45], char4[45]};
    char[174] <= {char44_0[46], char44_1[46], char44_2[46], char44_3[46], char44_4[46], char4[46]};
    char[175] <= {char44_0[47], char44_1[47], char44_2[47], char44_3[47], char44_4[47], char4[47]};
    char[176] <= {char44_0[48], char44_1[48], char44_2[48], char44_3[48], char44_4[48], char4[48]};
    char[177] <= {char44_0[49], char44_1[49], char44_2[49], char44_3[49], char44_4[49], char4[49]};
    char[178] <= {char44_0[50], char44_1[50], char44_2[50], char44_3[50], char44_4[50], char4[50]};
    char[179] <= {char44_0[51], char44_1[51], char44_2[51], char44_3[51], char44_4[51], char4[51]};
    char[180] <= {char44_0[52], char44_1[52], char44_2[52], char44_3[52], char44_4[52], char4[52]};
    char[181] <= {char44_0[53], char44_1[53], char44_2[53], char44_3[53], char44_4[53], char4[53]};
    char[182] <= {char44_0[54], char44_1[54], char44_2[54], char44_3[54], char44_4[54], char4[54]};
    char[183] <= {char44_0[55], char44_1[55], char44_2[55], char44_3[55], char44_4[55], char4[55]};
    char[184] <= {char44_0[56], char44_1[56], char44_2[56], char44_3[56], char44_4[56], char4[56]};
    char[185] <= {char44_0[57], char44_1[57], char44_2[57], char44_3[57], char44_4[57], char4[57]};
    char[186] <= {char44_0[58], char44_1[58], char44_2[58], char44_3[58], char44_4[58], char4[58]};
    char[187] <= {char44_0[59], char44_1[59], char44_2[59], char44_3[59], char44_4[59], char4[59]};
    char[188] <= {char44_0[60], char44_1[60], char44_2[60], char44_3[60], char44_4[60], char4[60]};
    char[189] <= {char44_0[61], char44_1[61], char44_2[61], char44_3[61], char44_4[61], char4[61]};
    char[190] <= {char44_0[62], char44_1[62], char44_2[62], char44_3[62], char44_4[62], char4[62]};
    char[191] <= {char44_0[63], char44_1[63], char44_2[63], char44_3[63], char44_4[63], char4[63]};


    char[192] <= 512'h0;
    char[193] <= 512'h0;
    char[194] <= 512'h0;
    char[195] <= 512'h0;
    char[196] <= 512'h0;
    char[197] <= 512'h0;
    char[198] <= 512'h0;
    char[199] <= 512'h0;
    char[200] <= 512'h0;
    char[201] <= 512'h0;
    char[202] <= 512'h0;
    char[203] <= 512'h0;
    char[204] <= 512'h0;
    char[205] <= 512'h0;
    char[206] <= 512'h0;
    char[207] <= 512'h0;
    char[208] <= 512'h0;
    char[209] <= 512'h0;
    char[210] <= 512'h0;
    char[211] <= 512'h0;
    char[212] <= 512'h0;
    char[213] <= 512'h0;
    char[214] <= 512'h0;
    char[215] <= 512'h0;
    char[216] <= 512'h0;
    char[217] <= 512'h0;
    char[218] <= 512'h0;
    char[219] <= 512'h0;
    char[220] <= 512'h0;
    char[221] <= 512'h0;
    char[222] <= 512'h0;
    char[223] <= 512'h0;
    char[224] <= 512'h0;
    char[225] <= 512'h0;
    char[226] <= 512'h0;
    char[227] <= 512'h0;
    char[228] <= 512'h0;
    char[229] <= 512'h0;
    char[230] <= 512'h0;
    char[231] <= 512'h0;
    char[232] <= 512'h0;
    char[233] <= 512'h0;
    char[234] <= 512'h0;
    char[235] <= 512'h0;
    char[236] <= 512'h0;
    char[237] <= 512'h0;
    char[238] <= 512'h0;
    char[239] <= 512'h0;
    char[240] <= 512'h0;
    char[241] <= 512'h0;
    char[242] <= 512'h0;
    char[243] <= 512'h0;
    char[244] <= 512'h0;
    char[245] <= 512'h0;
    char[246] <= 512'h0;
    char[247] <= 512'h0;
    char[248] <= 512'h0;
    char[249] <= 512'h0;
    char[250] <= 512'h0;
    char[251] <= 512'h0;
    char[252] <= 512'h0;
    char[253] <= 512'h0;
    char[254] <= 512'h0;
    char[255] <= 512'h0;
    char[256] <= 512'h0;
    char[257] <= 512'h0;
    char[258] <= 512'h0;
    char[259] <= 512'h0;
    char[260] <= 512'h0;
    char[261] <= 512'h0;
    char[262] <= 512'h0;
    char[263] <= 512'h0;
    char[264] <= 512'h0;
    char[265] <= 512'h0;
    char[266] <= 512'h0;
    char[267] <= 512'h0;
    char[268] <= 512'h0;
    char[269] <= 512'h0;
    char[270] <= 512'h0;
    char[271] <= 512'h0;
    char[272] <= 512'h0;
    char[273] <= 512'h0;
    char[274] <= 512'h0;
    char[275] <= 512'h0;
    char[276] <= 512'h0;
    char[277] <= 512'h0;
    char[278] <= 512'h0;
    char[279] <= 512'h0;
    char[280] <= 512'h0;
    char[281] <= 512'h0;
    char[282] <= 512'h0;
    char[283] <= 512'h0;
    char[284] <= 512'h0;
    char[285] <= 512'h0;
    char[286] <= 512'h0;
    char[287] <= 512'h0;
    char[288] <= 512'h0;
    char[289] <= 512'h0;
    char[290] <= 512'h0;
    char[291] <= 512'h0;
    char[292] <= 512'h0;
    char[293] <= 512'h0;
    char[294] <= 512'h0;
    char[295] <= 512'h0;
    char[296] <= 512'h0;
    char[297] <= 512'h0;
    char[298] <= 512'h0;
    char[299] <= 512'h0;
    char[300] <= 512'h0;
    char[301] <= 512'h0;
    char[302] <= 512'h0;
    char[303] <= 512'h0;
    char[304] <= 512'h0;
    char[305] <= 512'h0;
    char[306] <= 512'h0;
    char[307] <= 512'h0;
    char[308] <= 512'h0;
    char[309] <= 512'h0;
    char[310] <= 512'h0;
    char[311] <= 512'h0;
    char[312] <= 512'h0;
    char[313] <= 512'h0;
    char[314] <= 512'h0;
    char[315] <= 512'h0;
    char[316] <= 512'h0;
    char[317] <= 512'h0;
    char[318] <= 512'h0;
    char[319] <= 512'h0;
     char[320] <= 512'h0;
     char[321] <= 512'h0;
     char[322] <= 512'h0;
     char[323] <= 512'h0;
     char[324] <= 512'h0;
     char[325] <= 512'h0;
     char[326] <= 512'h0;
     char[327] <= 512'h0;
     char[328] <= 512'h0;
     char[329] <= 512'h0;
     char[330] <= 512'h0;
     char[331] <= 512'h0;
     char[332] <= 512'h0;
     char[333] <= 512'h0;
     char[334] <= 512'h0;
     char[335] <= 512'h0;
     char[336] <= 512'h0;
     char[337] <= 512'h0;
     char[338] <= 512'h0;
     char[339] <= 512'h0;
     char[340] <= 512'h0;
     char[341] <= 512'h0;
     char[342] <= 512'h0;
     char[343] <= 512'h0;
     char[344] <= 512'h0;
     char[345] <= 512'h0;
     char[346] <= 512'h0;
     char[347] <= 512'h0;
     char[348] <= 512'h0;
     char[349] <= 512'h0;
     char[350] <= 512'h0;
     char[351] <= 512'h0;
     char[352] <= 512'h0;
     char[353] <= 512'h0;
     char[354] <= 512'h0;
     char[355] <= 512'h0;
     char[356] <= 512'h0;
     char[357] <= 512'h0;
     char[358] <= 512'h0;
     char[359] <= 512'h0;
     char[360] <= 512'h0;
     char[361] <= 512'h0;
     char[362] <= 512'h0;
     char[363] <= 512'h0;
     char[364] <= 512'h0;
     char[365] <= 512'h0;
     char[366] <= 512'h0;
     char[367] <= 512'h0;
     char[368] <= 512'h0;
     char[369] <= 512'h0;
     char[370] <= 512'h0;
     char[371] <= 512'h0;
     char[372] <= 512'h0;
     char[373] <= 512'h0;
     char[374] <= 512'h0;
     char[375] <= 512'h0;
     char[376] <= 512'h0;
     char[377] <= 512'h0;
     char[378] <= 512'h0;
     char[379] <= 512'h0;
     char[380] <= 512'h0;
     char[381] <= 512'h0;
     char[382] <= 512'h0;
     char[383] <= 512'h0;
     char[384] <= 512'h0;
     char[385] <= 512'h0;
     char[386] <= 512'h0;
     char[387] <= 512'h0;
     char[388] <= 512'h0;
     char[389] <= 512'h0;
     char[390] <= 512'h0;
     char[391] <= 512'h0;
     char[392] <= 512'h0;
     char[393] <= 512'h0;
     char[394] <= 512'h0;
     char[395] <= 512'h0;
     char[396] <= 512'h0;
     char[397] <= 512'h0;
     char[398] <= 512'h0;
     char[399] <= 512'h0;
     char[400] <= 512'h0;
     char[401] <= 512'h0;
     char[402] <= 512'h0;
     char[403] <= 512'h0;
     char[404] <= 512'h0;
     char[405] <= 512'h0;
     char[406] <= 512'h0;
     char[407] <= 512'h0;
     char[408] <= 512'h0;
     char[409] <= 512'h0;
     char[410] <= 512'h0;
     char[411] <= 512'h0;
     char[412] <= 512'h0;
     char[413] <= 512'h0;
     char[414] <= 512'h0;
     char[415] <= 512'h0;
     char[416] <= 512'h0;
     char[417] <= 512'h0;
     char[418] <= 512'h0;
     char[419] <= 512'h0;
     char[420] <= 512'h0;
     char[421] <= 512'h0;
     char[422] <= 512'h0;
     char[423] <= 512'h0;
     char[424] <= 512'h0;
     char[425] <= 512'h0;
     char[426] <= 512'h0;
     char[427] <= 512'h0;
     char[428] <= 512'h0;
     char[429] <= 512'h0;
     char[430] <= 512'h0;
     char[431] <= 512'h0;
     char[432] <= 512'h0;
     char[433] <= 512'h0;
     char[434] <= 512'h0;
     char[435] <= 512'h0;
     char[436] <= 512'h0;
     char[437] <= 512'h0;
     char[438] <= 512'h0;
     char[439] <= 512'h0;
     char[440] <= 512'h0;
     char[441] <= 512'h0;
     char[442] <= 512'h0;
     char[443] <= 512'h0;
     char[444] <= 512'h0;
     char[445] <= 512'h0;
     char[446] <= 512'h0;
     char[447] <= 512'h0;
     char[448] <= 512'h0;
     char[449] <= 512'h0;
     char[450] <= 512'h0;
     char[451] <= 512'h0;
     char[452] <= 512'h0;
     char[453] <= 512'h0;
     char[454] <= 512'h0;
     char[455] <= 512'h0;
     char[456] <= 512'h0;
     char[457] <= 512'h0;
     char[458] <= 512'h0;
     char[459] <= 512'h0;
     char[460] <= 512'h0;
     char[461] <= 512'h0;
     char[462] <= 512'h0;
     char[463] <= 512'h0;
     char[464] <= 512'h0;
     char[465] <= 512'h0;
     char[466] <= 512'h0;
     char[467] <= 512'h0;
     char[468] <= 512'h0;
     char[469] <= 512'h0;
     char[470] <= 512'h0;
     char[471] <= 512'h0;
     char[472] <= 512'h0;
     char[473] <= 512'h0;
     char[474] <= 512'h0;
     char[475] <= 512'h0;
     char[476] <= 512'h0;
     char[477] <= 512'h0;
     char[478] <= 512'h0;
     char[479] <= 512'h0;
     
 
end

always @(posedge vga_clk , posedge sys_rst) begin
     if(sys_rst)begin
        pix_data <=black;
     end
     else if (pix_x<512 && char[pix_y][10'd255-pix_x] == 1'b1)
        /*if (pix_x >=416 && pix_y >= 128) pix_data <= white;
        else */pix_data <=blue;
     else
        pix_data <=white;
     
        
end

endmodule

module vga(//clk ��25MHZ
input wire sys_clk,//10oMhzʱ��
input wire sys_rst,//reset

input [31:0] a0,
input [31:0] a1,
input [31:0] a2,

output wire hsync,
output wire vsync,
output wire [11:0]vga_rgb
);
wire [9:0] pix_x;
wire [9:0] pix_y;
wire [11:0] pix_data;
wire clk_25m;

vga_control vc(
clk_25m ,  sys_rst ,  pix_data  ,  pix_x  , pix_y  , hsync,  vsync  ,  vga_rgb   
);

vga_draw vd(
clk_25m , sys_rst , a0, a1, a2  ,  pix_x , pix_y , pix_data
 );
 
Get25Clk Gc(
sys_clk  ,sys_rst ,clk_25m
);

endmodule

module Get25Clk(input sys_clk,input rst,output reg clk_25m);//��Ƶ��

parameter period =4;
reg[3:0] cnt;
always@(posedge sys_clk,posedge rst )begin
    if(rst)begin
        cnt<=0;
        clk_25m<=0;
        end
     else
           if(cnt==((period>>1)-1)) begin
           clk_25m <=~clk_25m;
           cnt<= 0;
           end 
           else begin
            cnt<=cnt+1;
            end
     end
endmodule
